<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>328.298,-195.234,402.227,-240.8</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>361.5,-196</position>
<gparam>LABEL_TEXT Circuits with Feedback</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_INVERTER</type>
<position>358,-208</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_INVERTER</type>
<position>372,-208</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>381,-208</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>345,-208</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>HE_JUNC_4</type>
<position>377,-208</position>
<input>
<ID>N_in0</ID>9 </input>
<input>
<ID>N_in1</ID>10 </input>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>HE_JUNC_4</type>
<position>354,-208</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>11 </input>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>358,-217.5</position>
<gparam>LABEL_TEXT Stable Feedback Circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>339,-232</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>391.5,-232</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_INVERTER</type>
<position>353,-232</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_INVERTER</type>
<position>366.5,-232</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_INVERTER</type>
<position>379,-232</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>HE_JUNC_4</type>
<position>348,-232</position>
<input>
<ID>N_in0</ID>18 </input>
<input>
<ID>N_in1</ID>17 </input>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>HE_JUNC_4</type>
<position>384.5,-232</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>15 </input>
<input>
<ID>N_in3</ID>19 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>365.5,-239</position>
<gparam>LABEL_TEXT Unstable Feedback Circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361,-208,369,-208</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354,-202.5,377,-202.5</points>
<intersection>354 4</intersection>
<intersection>377 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>377,-207,377,-202.5</points>
<connection>
<GID>12</GID>
<name>N_in3</name></connection>
<intersection>-202.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>354,-207,354,-202.5</points>
<connection>
<GID>13</GID>
<name>N_in3</name></connection>
<intersection>-202.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>375,-208,376,-208</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>378,-208,380,-208</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>12</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>355,-208,355,-208</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>347,-208,353,-208</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>13</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>369.5,-232,376,-232</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>356,-232,363.5,-232</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>385.5,-232,390.5,-232</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>382,-232,383.5,-232</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>21</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,-232,350,-232</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>341,-232,347,-232</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>348,-227.5,384.5,-227.5</points>
<intersection>348 4</intersection>
<intersection>384.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>384.5,-231,384.5,-227.5</points>
<connection>
<GID>21</GID>
<name>N_in3</name></connection>
<intersection>-227.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>348,-231,348,-227.5</points>
<connection>
<GID>20</GID>
<name>N_in3</name></connection>
<intersection>-227.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>124.226,-40.9918,196.317,-85.425</PageViewport>
<gate>
<ID>386</ID>
<type>AA_LABEL</type>
<position>164.5,-61.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>842</ID>
<type>AA_LABEL</type>
<position>138,-71.5</position>
<gparam>LABEL_TEXT S=0,R=0 not allowed</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>144,-44.5</position>
<gparam>LABEL_TEXT Quiescent state R=1 S=1 (holds value of Q)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>142.5,-67.5</position>
<gparam>LABEL_TEXT Set S=0 (R=1) and reset back to S=1 </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>143.5,-47</position>
<gparam>LABEL_TEXT Set R=0, S=1 and reset back to R=1 ??</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>BA_NAND2</type>
<position>148,-54</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>BA_NAND2</type>
<position>148.5,-62</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>HA_JUNC_2</type>
<position>140.5,-53</position>
<input>
<ID>N_in0</ID>83 </input>
<input>
<ID>N_in1</ID>76 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>HA_JUNC_2</type>
<position>140.5,-63</position>
<input>
<ID>N_in0</ID>82 </input>
<input>
<ID>N_in1</ID>77 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>HE_JUNC_4</type>
<position>153,-62</position>
<input>
<ID>N_in0</ID>78 </input>
<input>
<ID>N_in1</ID>290 </input>
<input>
<ID>N_in3</ID>79 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>HE_JUNC_4</type>
<position>153.5,-54</position>
<input>
<ID>N_in0</ID>80 </input>
<input>
<ID>N_in1</ID>84 </input>
<input>
<ID>N_in2</ID>81 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>134.5,-53</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>135.5,-63</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>159.5,-54</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>132.5,-53</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>133,-63</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>144.5,-41.5</position>
<gparam>LABEL_TEXT RS  Latch</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>379</ID>
<type>GA_LED</type>
<position>159.5,-62</position>
<input>
<ID>N_in0</ID>290 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>384</ID>
<type>AA_LABEL</type>
<position>163.5,-53.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-53,145,-53</points>
<connection>
<GID>104</GID>
<name>N_in1</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>141.5,-63,145.5,-63</points>
<connection>
<GID>105</GID>
<name>N_in1</name></connection>
<connection>
<GID>103</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151.5,-62,152,-62</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-61,153,-57.5</points>
<connection>
<GID>106</GID>
<name>N_in3</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-57.5,153,-57.5</points>
<intersection>145 2</intersection>
<intersection>153 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>145,-57.5,145,-55</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>-57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>151,-54,152.5,-54</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>107</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-61,143,-56.5</points>
<intersection>-61 1</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-61,145.5,-61</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-56.5,153.5,-56.5</points>
<intersection>143 0</intersection>
<intersection>153.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>153.5,-56.5,153.5,-55</points>
<connection>
<GID>107</GID>
<name>N_in2</name></connection>
<intersection>-56.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-63,139.5,-63</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<connection>
<GID>105</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136.5,-53,139.5,-53</points>
<connection>
<GID>104</GID>
<name>N_in0</name></connection>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154.5,-54,158.5,-54</points>
<connection>
<GID>107</GID>
<name>N_in1</name></connection>
<connection>
<GID>111</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-62,158.5,-62</points>
<connection>
<GID>379</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>N_in1</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-61,-2.75657,16.1,-50.277</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-39.5,-22.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>-30,-30.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>-6,-21.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>-4,-34</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>-1,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>BA_NAND2</type>
<position>-0.5,-32</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>HA_JUNC_2</type>
<position>-8.5,-23</position>
<input>
<ID>N_in0</ID>45 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>HA_JUNC_2</type>
<position>-8.5,-33</position>
<input>
<ID>N_in0</ID>46 </input>
<input>
<ID>N_in1</ID>5 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>HE_JUNC_4</type>
<position>4,-32</position>
<input>
<ID>N_in0</ID>6 </input>
<input>
<ID>N_in3</ID>20 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>HE_JUNC_4</type>
<position>4.5,-24</position>
<input>
<ID>N_in0</ID>37 </input>
<input>
<ID>N_in1</ID>39 </input>
<input>
<ID>N_in2</ID>38 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>10.5,-24</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-40,-19</position>
<gparam>LABEL_TEXT D  (input)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>BA_NAND2</type>
<position>-18.5,-23.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>BA_NAND2</type>
<position>-18.5,-33.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_SMALL_INVERTER</type>
<position>-24,-34.5</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>HE_JUNC_4</type>
<position>-26,-22.5</position>
<input>
<ID>N_in0</ID>3 </input>
<input>
<ID>N_in1</ID>41 </input>
<input>
<ID>N_in2</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>HE_JUNC_4</type>
<position>-22,-28.5</position>
<input>
<ID>N_in0</ID>47 </input>
<input>
<ID>N_in2</ID>44 </input>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>-46,-28.5</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>-51,-34.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>-14,-12</position>
<gparam>LABEL_TEXT D Latch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>11.5,-20.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>-16.5,-40</position>
<gparam>LABEL_TEXT Value of Q = value of D stored when WE=1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-22.5,-27,-22.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7.5,-23,-4,-23</points>
<connection>
<GID>23</GID>
<name>N_in1</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7.5,-33,-3.5,-33</points>
<connection>
<GID>24</GID>
<name>N_in1</name></connection>
<connection>
<GID>7</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>2.5,-32,3,-32</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<connection>
<GID>25</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-31,4,-27.5</points>
<connection>
<GID>25</GID>
<name>N_in3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-27.5,4,-27.5</points>
<intersection>-4 2</intersection>
<intersection>4 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-4,-27.5,-4,-25</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>2,-24,3.5,-24</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-31,-6,-26.5</points>
<intersection>-31 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-31,-3.5,-31</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6,-26.5,4.5,-26.5</points>
<intersection>-6 0</intersection>
<intersection>4.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-26.5,4.5,-25</points>
<connection>
<GID>26</GID>
<name>N_in2</name></connection>
<intersection>-26.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>5.5,-24,9.5,-24</points>
<connection>
<GID>26</GID>
<name>N_in1</name></connection>
<connection>
<GID>27</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-22,-34.5,-21.5,-34.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-25,-22.5,-21.5,-22.5</points>
<connection>
<GID>32</GID>
<name>N_in1</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-34.5,-26,-23.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-27.5,-22,-24.5</points>
<connection>
<GID>55</GID>
<name>N_in3</name></connection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-24.5,-21.5,-24.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-32.5,-22,-29.5</points>
<connection>
<GID>55</GID>
<name>N_in2</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,-32.5,-21.5,-32.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-23.5,-12.5,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-23,-9.5,-23</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-23.5,-12.5,-23.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-33.5,-12.5,-33</points>
<intersection>-33.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-33,-9.5,-33</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15.5,-33.5,-12.5,-33.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-28.5,-23,-28.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>55</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>21.9489,0.02469,217.901,-120.75</PageViewport>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>124,-17.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>126,-30</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>BA_NAND2</type>
<position>129,-20</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>BA_NAND2</type>
<position>129.5,-28</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>HA_JUNC_2</type>
<position>121.5,-19</position>
<input>
<ID>N_in0</ID>130 </input>
<input>
<ID>N_in1</ID>118 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>HA_JUNC_2</type>
<position>121.5,-29</position>
<input>
<ID>N_in0</ID>131 </input>
<input>
<ID>N_in1</ID>119 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>HE_JUNC_4</type>
<position>134,-28</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in3</ID>121 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>HE_JUNC_4</type>
<position>134.5,-20</position>
<input>
<ID>N_in0</ID>122 </input>
<input>
<ID>N_in1</ID>124 </input>
<input>
<ID>N_in2</ID>123 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>140.5,-20</position>
<input>
<ID>N_in0</ID>124 </input>
<input>
<ID>N_in1</ID>140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>104,-15.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>111.5,-19.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>BA_NAND2</type>
<position>111.5,-29.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>125 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_SMALL_INVERTER</type>
<position>106,-30.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>75</ID>
<type>HE_JUNC_4</type>
<position>106,-18.5</position>
<input>
<ID>N_in0</ID>133 </input>
<input>
<ID>N_in1</ID>126 </input>
<input>
<ID>N_in2</ID>127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>HE_JUNC_4</type>
<position>108,-24.5</position>
<input>
<ID>N_in0</ID>132 </input>
<input>
<ID>N_in2</ID>129 </input>
<input>
<ID>N_in3</ID>128 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>DD_KEYPAD_HEX</type>
<position>66,-55</position>
<output>
<ID>OUT_0</ID>136 </output>
<output>
<ID>OUT_1</ID>135 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>133 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 12</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>86,-119.5</position>
<output>
<ID>OUT_0</ID>132 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>85</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>180,-54.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>140 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 12</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>100.5,-49.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>124.5,-40.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>126.5,-53</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>BA_NAND2</type>
<position>129.5,-43</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>124,-1</position>
<gparam>LABEL_TEXT 4 bit register using D latches</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>BA_NAND2</type>
<position>130,-51</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>HA_JUNC_2</type>
<position>122,-42</position>
<input>
<ID>N_in0</ID>75 </input>
<input>
<ID>N_in1</ID>48 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>122,-52</position>
<input>
<ID>N_in0</ID>85 </input>
<input>
<ID>N_in1</ID>49 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>HE_JUNC_4</type>
<position>134.5,-51</position>
<input>
<ID>N_in0</ID>50 </input>
<input>
<ID>N_in3</ID>51 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>HE_JUNC_4</type>
<position>135,-43</position>
<input>
<ID>N_in0</ID>52 </input>
<input>
<ID>N_in1</ID>66 </input>
<input>
<ID>N_in2</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>141,-43</position>
<input>
<ID>N_in0</ID>66 </input>
<input>
<ID>N_in1</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>BA_NAND2</type>
<position>112,-42.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_NAND2</type>
<position>112,-52.5</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>106.5,-53.5</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>HE_JUNC_4</type>
<position>106.5,-41.5</position>
<input>
<ID>N_in0</ID>134 </input>
<input>
<ID>N_in1</ID>71 </input>
<input>
<ID>N_in2</ID>72 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>HE_JUNC_4</type>
<position>108.5,-47.5</position>
<input>
<ID>N_in0</ID>132 </input>
<input>
<ID>N_in2</ID>74 </input>
<input>
<ID>N_in3</ID>73 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>100,-72.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>63.5,-44</position>
<gparam>LABEL_TEXT Keypad</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>124,-63.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>126,-76</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AA_LABEL</type>
<position>73.5,-117</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>BA_NAND2</type>
<position>129,-66</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>BA_NAND2</type>
<position>129.5,-74</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>HA_JUNC_2</type>
<position>121.5,-65</position>
<input>
<ID>N_in0</ID>102 </input>
<input>
<ID>N_in1</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>HA_JUNC_2</type>
<position>121.5,-75</position>
<input>
<ID>N_in0</ID>103 </input>
<input>
<ID>N_in1</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>HE_JUNC_4</type>
<position>134,-74</position>
<input>
<ID>N_in0</ID>92 </input>
<input>
<ID>N_in3</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>HE_JUNC_4</type>
<position>134.5,-66</position>
<input>
<ID>N_in0</ID>94 </input>
<input>
<ID>N_in1</ID>96 </input>
<input>
<ID>N_in2</ID>95 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>140.5,-66</position>
<input>
<ID>N_in0</ID>96 </input>
<input>
<ID>N_in1</ID>138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>AA_LABEL</type>
<position>101,-64.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>BA_NAND2</type>
<position>111.5,-65.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>BA_NAND2</type>
<position>111.5,-76.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AE_SMALL_INVERTER</type>
<position>106,-76.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>154</ID>
<type>HE_JUNC_4</type>
<position>106,-64.5</position>
<input>
<ID>N_in0</ID>135 </input>
<input>
<ID>N_in1</ID>98 </input>
<input>
<ID>N_in2</ID>99 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>HE_JUNC_4</type>
<position>108,-70.5</position>
<input>
<ID>N_in0</ID>132 </input>
<input>
<ID>N_in2</ID>101 </input>
<input>
<ID>N_in3</ID>100 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>102,-94</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>126,-85</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>128,-97.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>116,-8</position>
<gparam>LABEL_TEXT D Latch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>BA_NAND2</type>
<position>131,-87.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>BA_NAND2</type>
<position>131.5,-95.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>HA_JUNC_2</type>
<position>123.5,-86.5</position>
<input>
<ID>N_in0</ID>116 </input>
<input>
<ID>N_in1</ID>104 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>HA_JUNC_2</type>
<position>123.5,-96.5</position>
<input>
<ID>N_in0</ID>117 </input>
<input>
<ID>N_in1</ID>105 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>HE_JUNC_4</type>
<position>136,-95.5</position>
<input>
<ID>N_in0</ID>106 </input>
<input>
<ID>N_in3</ID>107 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>HE_JUNC_4</type>
<position>136.5,-87.5</position>
<input>
<ID>N_in0</ID>108 </input>
<input>
<ID>N_in1</ID>110 </input>
<input>
<ID>N_in2</ID>109 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>142.5,-87.5</position>
<input>
<ID>N_in0</ID>110 </input>
<input>
<ID>N_in1</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>103,-86</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>BA_NAND2</type>
<position>113.5,-87</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>BA_NAND2</type>
<position>113.5,-97</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AE_SMALL_INVERTER</type>
<position>108,-98</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>171</ID>
<type>HE_JUNC_4</type>
<position>108,-86</position>
<input>
<ID>N_in0</ID>136 </input>
<input>
<ID>N_in1</ID>112 </input>
<input>
<ID>N_in2</ID>113 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>HE_JUNC_4</type>
<position>110,-92</position>
<input>
<ID>N_in0</ID>132 </input>
<input>
<ID>N_in2</ID>115 </input>
<input>
<ID>N_in3</ID>114 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>100,-26.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-42,126.5,-42</points>
<connection>
<GID>126</GID>
<name>N_in1</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123,-52,127,-52</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<connection>
<GID>125</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>133,-51,133.5,-51</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-50,134.5,-46.5</points>
<connection>
<GID>128</GID>
<name>N_in3</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,-46.5,134.5,-46.5</points>
<intersection>126.5 2</intersection>
<intersection>134.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126.5,-46.5,126.5,-44</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132.5,-43,134,-43</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-50,124.5,-45.5</points>
<intersection>-50 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-50,127,-50</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-45.5,135,-45.5</points>
<intersection>124.5 0</intersection>
<intersection>135 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>135,-45.5,135,-44</points>
<connection>
<GID>129</GID>
<name>N_in2</name></connection>
<intersection>-45.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>136,-43,140,-43</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<connection>
<GID>131</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-53.5,109,-53.5</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107.5,-41.5,109,-41.5</points>
<connection>
<GID>136</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-53.5,104.5,-42.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-42.5,106.5,-42.5</points>
<connection>
<GID>136</GID>
<name>N_in2</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-46.5,108.5,-43.5</points>
<connection>
<GID>137</GID>
<name>N_in3</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-43.5,109,-43.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-51.5,108.5,-48.5</points>
<connection>
<GID>137</GID>
<name>N_in2</name></connection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-51.5,109,-51.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-42.5,118,-42</points>
<intersection>-42.5 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-42,121,-42</points>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-42.5,118,-42.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-52.5,118,-52</points>
<intersection>-52.5 2</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-52,121,-52</points>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,-52.5,118,-52.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-65,126,-65</points>
<connection>
<GID>145</GID>
<name>N_in1</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-75,126.5,-75</points>
<connection>
<GID>146</GID>
<name>N_in1</name></connection>
<connection>
<GID>144</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132.5,-74,133,-74</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>147</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-73,134,-69.5</points>
<connection>
<GID>147</GID>
<name>N_in3</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-69.5,134,-69.5</points>
<intersection>126 2</intersection>
<intersection>134 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-69.5,126,-67</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>-69.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132,-66,133.5,-66</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-73,124,-68.5</points>
<intersection>-73 1</intersection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-73,126.5,-73</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124,-68.5,134.5,-68.5</points>
<intersection>124 0</intersection>
<intersection>134.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-68.5,134.5,-67</points>
<connection>
<GID>148</GID>
<name>N_in2</name></connection>
<intersection>-68.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>135.5,-66,139.5,-66</points>
<connection>
<GID>148</GID>
<name>N_in1</name></connection>
<connection>
<GID>149</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-77.5,108.5,-77.5</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,-77.5,108,-76.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>107,-64.5,108.5,-64.5</points>
<connection>
<GID>154</GID>
<name>N_in1</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-76.5,104,-65.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-65.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,-65.5,106,-65.5</points>
<connection>
<GID>154</GID>
<name>N_in2</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-69.5,108,-66.5</points>
<connection>
<GID>155</GID>
<name>N_in3</name></connection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-66.5,108.5,-66.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-75.5,108,-71.5</points>
<connection>
<GID>155</GID>
<name>N_in2</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-75.5,108.5,-75.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-65.5,117.5,-65</points>
<intersection>-65.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-65,120.5,-65</points>
<connection>
<GID>145</GID>
<name>N_in0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-65.5,117.5,-65.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-76.5,117.5,-75</points>
<intersection>-76.5 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-75,120.5,-75</points>
<connection>
<GID>146</GID>
<name>N_in0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-76.5,117.5,-76.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-86.5,128,-86.5</points>
<connection>
<GID>162</GID>
<name>N_in1</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-96.5,128.5,-96.5</points>
<connection>
<GID>163</GID>
<name>N_in1</name></connection>
<connection>
<GID>161</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>134.5,-95.5,135,-95.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<connection>
<GID>164</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-97.5,136,-94.5</points>
<connection>
<GID>164</GID>
<name>N_in3</name></connection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-97.5,136,-97.5</points>
<intersection>127 2</intersection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>127,-97.5,127,-88.5</points>
<intersection>-97.5 1</intersection>
<intersection>-88.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>127,-88.5,128,-88.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>127 2</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>134,-87.5,135.5,-87.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-96.5,125,-94.5</points>
<intersection>-96.5 2</intersection>
<intersection>-94.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-94.5,128.5,-94.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-96.5,136.5,-96.5</points>
<intersection>125 0</intersection>
<intersection>136.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>136.5,-96.5,136.5,-88.5</points>
<connection>
<GID>165</GID>
<name>N_in2</name></connection>
<intersection>-96.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>137.5,-87.5,141.5,-87.5</points>
<connection>
<GID>165</GID>
<name>N_in1</name></connection>
<connection>
<GID>166</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>110,-98,110.5,-98</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<connection>
<GID>169</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-86,110.5,-86</points>
<connection>
<GID>171</GID>
<name>N_in1</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-98,106,-87</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>106,-87,108,-87</points>
<connection>
<GID>171</GID>
<name>N_in2</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-91,110,-88</points>
<connection>
<GID>172</GID>
<name>N_in3</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-88,110.5,-88</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-96,110,-93</points>
<connection>
<GID>172</GID>
<name>N_in2</name></connection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-96,110.5,-96</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>110 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-87,119.5,-86.5</points>
<intersection>-87 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-86.5,122.5,-86.5</points>
<connection>
<GID>162</GID>
<name>N_in0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-87,119.5,-87</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-97,119.5,-96.5</points>
<intersection>-97 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-96.5,122.5,-96.5</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<intersection>119.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-97,119.5,-97</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-19,126,-19</points>
<connection>
<GID>66</GID>
<name>N_in1</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-29,126.5,-29</points>
<connection>
<GID>67</GID>
<name>N_in1</name></connection>
<connection>
<GID>65</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132.5,-28,133,-28</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-27,134,-23.5</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-23.5,134,-23.5</points>
<intersection>126 2</intersection>
<intersection>134 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126,-23.5,126,-21</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>132,-20,133.5,-20</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-27,124,-22.5</points>
<intersection>-27 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-27,126.5,-27</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124,-22.5,134.5,-22.5</points>
<intersection>124 0</intersection>
<intersection>134.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-22.5,134.5,-21</points>
<connection>
<GID>69</GID>
<name>N_in2</name></connection>
<intersection>-22.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>135.5,-20,139.5,-20</points>
<connection>
<GID>69</GID>
<name>N_in1</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108,-30.5,108.5,-30.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>107,-18.5,108.5,-18.5</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<connection>
<GID>72</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-30.5,104,-19.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,-19.5,106,-19.5</points>
<connection>
<GID>75</GID>
<name>N_in2</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-23.5,108,-20.5</points>
<connection>
<GID>76</GID>
<name>N_in3</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-20.5,108.5,-20.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-28.5,108,-25.5</points>
<connection>
<GID>76</GID>
<name>N_in2</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-28.5,108.5,-28.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-19.5,117.5,-19</points>
<intersection>-19.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-19,120.5,-19</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-19.5,117.5,-19.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-29.5,117.5,-29</points>
<intersection>-29.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-29,120.5,-29</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-29.5,117.5,-29.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-119.5,97.5,-24.5</points>
<intersection>-119.5 1</intersection>
<intersection>-92 2</intersection>
<intersection>-70.5 4</intersection>
<intersection>-47.5 6</intersection>
<intersection>-24.5 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-119.5,97.5,-119.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-92,109,-92</points>
<connection>
<GID>172</GID>
<name>N_in0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>97.5,-70.5,107,-70.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>97.5,-47.5,107.5,-47.5</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>97.5,-24.5,107,-24.5</points>
<connection>
<GID>76</GID>
<name>N_in0</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-52,79.5,-18.5</points>
<intersection>-52 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-18.5,105,-18.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-52,79.5,-52</points>
<connection>
<GID>77</GID>
<name>OUT_3</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-54,87.5,-41.5</points>
<intersection>-54 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-54,87.5,-54</points>
<connection>
<GID>77</GID>
<name>OUT_2</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-41.5,105.5,-41.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-64.5,87.5,-56</points>
<intersection>-64.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-56,87.5,-56</points>
<connection>
<GID>77</GID>
<name>OUT_1</name></connection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-64.5,105,-64.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-86,79.5,-58</points>
<intersection>-86 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-58,79.5,-58</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79.5,-86,107,-86</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>143.5,-87.5,177,-87.5</points>
<connection>
<GID>166</GID>
<name>N_in1</name></connection>
<intersection>177 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>177,-87.5,177,-55.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-87.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-66,173,-54.5</points>
<intersection>-66 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-66,173,-66</points>
<connection>
<GID>149</GID>
<name>N_in1</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>173,-54.5,177,-54.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-53.5,172.5,-43</points>
<intersection>-53.5 2</intersection>
<intersection>-43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-43,172.5,-43</points>
<connection>
<GID>131</GID>
<name>N_in1</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>172.5,-53.5,177,-53.5</points>
<connection>
<GID>85</GID>
<name>IN_2</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176.5,-52.5,176.5,-20</points>
<intersection>-52.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-20,176.5,-20</points>
<connection>
<GID>70</GID>
<name>N_in1</name></connection>
<intersection>176.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176.5,-52.5,177,-52.5</points>
<connection>
<GID>85</GID>
<name>IN_3</name></connection>
<intersection>176.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>56.284,-73.9753,358.69,-260.362</PageViewport>
<gate>
<ID>193</ID>
<type>BA_NAND2</type>
<position>179,-142</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>BA_NAND2</type>
<position>179,-152</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_SMALL_INVERTER</type>
<position>173.5,-153</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>HE_JUNC_4</type>
<position>171,-141</position>
<input>
<ID>N_in1</ID>151 </input>
<input>
<ID>N_in2</ID>152 </input>
<input>
<ID>N_in3</ID>142 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>HE_JUNC_4</type>
<position>175.5,-147</position>
<input>
<ID>N_in0</ID>209 </input>
<input>
<ID>N_in2</ID>154 </input>
<input>
<ID>N_in3</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>166.5,-174</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>191,-163</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>193,-175.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>BA_NAND2</type>
<position>196,-165.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>BA_NAND2</type>
<position>196.5,-173.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>HA_JUNC_2</type>
<position>188.5,-164.5</position>
<input>
<ID>N_in0</ID>168 </input>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>HA_JUNC_2</type>
<position>188.5,-174.5</position>
<input>
<ID>N_in0</ID>169 </input>
<input>
<ID>N_in1</ID>158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>HE_JUNC_4</type>
<position>201,-173.5</position>
<input>
<ID>N_in0</ID>159 </input>
<input>
<ID>N_in3</ID>160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>HE_JUNC_4</type>
<position>201.5,-165.5</position>
<input>
<ID>N_in0</ID>161 </input>
<input>
<ID>N_in1</ID>163 </input>
<input>
<ID>N_in2</ID>162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>207.5,-165.5</position>
<input>
<ID>N_in0</ID>163 </input>
<input>
<ID>N_in1</ID>211 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>168,-164</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>172,-95.5</position>
<gparam>LABEL_TEXT Memory: 4 locations, 1 bit addressability</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>BA_NAND2</type>
<position>178.5,-165</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>BA_NAND2</type>
<position>178.5,-176</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>137.5,-150</position>
<gparam>LABEL_TEXT Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AE_SMALL_INVERTER</type>
<position>173,-176</position>
<input>
<ID>IN_0</ID>200 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>HE_JUNC_4</type>
<position>171,-164</position>
<input>
<ID>N_in1</ID>165 </input>
<input>
<ID>N_in2</ID>200 </input>
<input>
<ID>N_in3</ID>152 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>HE_JUNC_4</type>
<position>175,-170</position>
<input>
<ID>N_in0</ID>201 </input>
<input>
<ID>N_in2</ID>167 </input>
<input>
<ID>N_in3</ID>166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>178.5,-191.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>193,-184.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>195,-197</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>183,-107.5</position>
<gparam>LABEL_TEXT D Latch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>BA_NAND2</type>
<position>198,-187</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>BA_NAND2</type>
<position>198.5,-195</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>HA_JUNC_2</type>
<position>190.5,-186</position>
<input>
<ID>N_in0</ID>182 </input>
<input>
<ID>N_in1</ID>170 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>HA_JUNC_2</type>
<position>190.5,-196</position>
<input>
<ID>N_in0</ID>183 </input>
<input>
<ID>N_in1</ID>171 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>HE_JUNC_4</type>
<position>203,-195</position>
<input>
<ID>N_in0</ID>172 </input>
<input>
<ID>N_in3</ID>173 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>HE_JUNC_4</type>
<position>203.5,-187</position>
<input>
<ID>N_in0</ID>174 </input>
<input>
<ID>N_in1</ID>176 </input>
<input>
<ID>N_in2</ID>175 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>GA_LED</type>
<position>209.5,-187</position>
<input>
<ID>N_in0</ID>176 </input>
<input>
<ID>N_in1</ID>210 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>168.5,-185</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>BA_NAND2</type>
<position>180.5,-186.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>BA_NAND2</type>
<position>180.5,-196.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-197.5</position>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>HE_JUNC_4</type>
<position>171,-185.5</position>
<input>
<ID>N_in1</ID>178 </input>
<input>
<ID>N_in2</ID>179 </input>
<input>
<ID>N_in3</ID>200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>HE_JUNC_4</type>
<position>177,-191.5</position>
<input>
<ID>N_in0</ID>202 </input>
<input>
<ID>N_in2</ID>181 </input>
<input>
<ID>N_in3</ID>180 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>177.5,-124</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>191,-117</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>193,-129.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>BA_NAND2</type>
<position>196,-119.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>BA_NAND2</type>
<position>196.5,-127.5</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>HA_JUNC_2</type>
<position>188.5,-118.5</position>
<input>
<ID>N_in0</ID>195 </input>
<input>
<ID>N_in1</ID>184 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AA_LABEL</type>
<position>171.5,-100.5</position>
<gparam>LABEL_TEXT each D-latch stores 1 bit at 1 location</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>HA_JUNC_2</type>
<position>188.5,-128.5</position>
<input>
<ID>N_in0</ID>196 </input>
<input>
<ID>N_in1</ID>185 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>HE_JUNC_4</type>
<position>201,-127.5</position>
<input>
<ID>N_in0</ID>186 </input>
<input>
<ID>N_in3</ID>187 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>HE_JUNC_4</type>
<position>201.5,-119.5</position>
<input>
<ID>N_in0</ID>188 </input>
<input>
<ID>N_in1</ID>190 </input>
<input>
<ID>N_in2</ID>189 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>GA_LED</type>
<position>207.5,-119.5</position>
<input>
<ID>N_in0</ID>190 </input>
<input>
<ID>N_in1</ID>213 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>171,-115</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>BA_NAND2</type>
<position>178.5,-119</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>GA_LED</type>
<position>251,-153.5</position>
<input>
<ID>N_in0</ID>214 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>BA_DECODER_2x4</type>
<position>134.5,-157</position>
<input>
<ID>ENABLE</ID>199 </input>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT_0</ID>208 </output>
<output>
<ID>OUT_1</ID>207 </output>
<output>
<ID>OUT_2</ID>206 </output>
<output>
<ID>OUT_3</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>117,-161</position>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>117,-157</position>
<output>
<ID>OUT_0</ID>198 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_TOGGLE</type>
<position>118,-151</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_AND2</type>
<position>166.5,-124</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_AND2</type>
<position>167.5,-146.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_AND2</type>
<position>166.5,-170</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>168.5,-191.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>138.5,-219</position>
<gparam>LABEL_TEXT Write/Read</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AA_TOGGLE</type>
<position>116.5,-110</position>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>104,-109</position>
<gparam>LABEL_TEXT Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>104,-112</position>
<gparam>LABEL_TEXT (to store)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AE_MUX_4x1</type>
<position>233.5,-153.5</position>
<input>
<ID>IN_0</ID>210 </input>
<input>
<ID>IN_1</ID>211 </input>
<input>
<ID>IN_2</ID>212 </input>
<input>
<ID>IN_3</ID>213 </input>
<output>
<ID>OUT</ID>214 </output>
<input>
<ID>SEL_0</ID>197 </input>
<input>
<ID>SEL_1</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>99,-156</position>
<gparam>LABEL_TEXT Memory Address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>236,-143.5</position>
<gparam>LABEL_TEXT Address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>BA_NAND2</type>
<position>178.5,-129</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>191 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_SMALL_INVERTER</type>
<position>173,-130</position>
<input>
<ID>IN_0</ID>142 </input>
<output>
<ID>OUT_0</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>HE_JUNC_4</type>
<position>171,-118</position>
<input>
<ID>N_in0</ID>205 </input>
<input>
<ID>N_in1</ID>192 </input>
<input>
<ID>N_in2</ID>142 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>HE_JUNC_4</type>
<position>175,-124</position>
<input>
<ID>N_in0</ID>141 </input>
<input>
<ID>N_in2</ID>194 </input>
<input>
<ID>N_in3</ID>193 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_TOGGLE</type>
<position>153,-219</position>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>167.5,-149</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>191.5,-140</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>193.5,-152.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>BA_NAND2</type>
<position>196.5,-142.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>BA_NAND2</type>
<position>197,-150.5</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>HA_JUNC_2</type>
<position>189,-141.5</position>
<input>
<ID>N_in0</ID>155 </input>
<input>
<ID>N_in1</ID>143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>HA_JUNC_2</type>
<position>189,-151.5</position>
<input>
<ID>N_in0</ID>156 </input>
<input>
<ID>N_in1</ID>144 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>HE_JUNC_4</type>
<position>201.5,-150.5</position>
<input>
<ID>N_in0</ID>145 </input>
<input>
<ID>N_in3</ID>146 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>HE_JUNC_4</type>
<position>202,-142.5</position>
<input>
<ID>N_in0</ID>147 </input>
<input>
<ID>N_in1</ID>149 </input>
<input>
<ID>N_in2</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>208,-142.5</position>
<input>
<ID>N_in0</ID>149 </input>
<input>
<ID>N_in1</ID>212 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-123,175,-120</points>
<connection>
<GID>181</GID>
<name>N_in3</name></connection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-120,175.5,-120</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-128,175,-125</points>
<connection>
<GID>181</GID>
<name>N_in2</name></connection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-128,175.5,-128</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-119,184.5,-118.5</points>
<intersection>-119 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-118.5,187.5,-118.5</points>
<connection>
<GID>238</GID>
<name>N_in0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-119,184.5,-119</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-129,184.5,-128.5</points>
<intersection>-129 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-128.5,187.5,-128.5</points>
<connection>
<GID>240</GID>
<name>N_in0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-129,184.5,-129</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-208,125,-161</points>
<intersection>-208 1</intersection>
<intersection>-161 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-208,240,-208</points>
<intersection>125 0</intersection>
<intersection>129 4</intersection>
<intersection>240 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-161,125,-161</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,-208,240,-148.5</points>
<intersection>-208 1</intersection>
<intersection>-148.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>129,-208,129,-158.5</points>
<intersection>-208 1</intersection>
<intersection>-158.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>234.5,-148.5,240,-148.5</points>
<connection>
<GID>175</GID>
<name>SEL_0</name></connection>
<intersection>240 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>129,-158.5,131.5,-158.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>129 4</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-211,121.5,-157</points>
<intersection>-211 1</intersection>
<intersection>-157 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-211,243.5,-211</points>
<intersection>121.5 0</intersection>
<intersection>131.5 4</intersection>
<intersection>243.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119,-157,121.5,-157</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>243.5,-211,243.5,-147</points>
<intersection>-211 1</intersection>
<intersection>-147 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>131.5,-211,131.5,-157.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>233.5,-147,243.5,-147</points>
<intersection>233.5 6</intersection>
<intersection>243.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>233.5,-148.5,233.5,-147</points>
<connection>
<GID>175</GID>
<name>SEL_1</name></connection>
<intersection>-147 5</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-155.5,125.5,-151</points>
<intersection>-155.5 1</intersection>
<intersection>-151 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125.5,-155.5,131.5,-155.5</points>
<connection>
<GID>247</GID>
<name>ENABLE</name></connection>
<intersection>125.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-151,125.5,-151</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-184.5,171,-165</points>
<connection>
<GID>231</GID>
<name>N_in3</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<connection>
<GID>214</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169.5,-170,174,-170</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<connection>
<GID>215</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>171.5,-191.5,176,-191.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159.5,-219,159.5,-125</points>
<intersection>-219 2</intersection>
<intersection>-192.5 5</intersection>
<intersection>-171 4</intersection>
<intersection>-147.5 3</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>159.5,-125,163.5,-125</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-219,159.5,-219</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>159.5,-147.5,164.5,-147.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>159.5,-171,163.5,-171</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<intersection>159.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>159.5,-192.5,165.5,-192.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>159.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-155.5,151,-123</points>
<intersection>-155.5 2</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-123,163.5,-123</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-155.5,151,-155.5</points>
<connection>
<GID>247</GID>
<name>OUT_3</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118.5,-110,171,-110</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>171 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>171,-118,171,-110</points>
<intersection>-118 4</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>170,-118,171,-118</points>
<connection>
<GID>180</GID>
<name>N_in0</name></connection>
<intersection>171 3</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152.5,-156.5,152.5,-145.5</points>
<intersection>-156.5 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152.5,-145.5,164.5,-145.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>152.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-156.5,152.5,-156.5</points>
<connection>
<GID>247</GID>
<name>OUT_2</name></connection>
<intersection>152.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>137.5,-157.5,163.5,-157.5</points>
<connection>
<GID>247</GID>
<name>OUT_1</name></connection>
<intersection>163.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>163.5,-169,163.5,-157.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,-190.5,151.5,-158.5</points>
<intersection>-190.5 2</intersection>
<intersection>-158.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-158.5,151.5,-158.5</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>151.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151.5,-190.5,165.5,-190.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>151.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172.5,-147,172.5,-146.5</points>
<intersection>-147 1</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>172.5,-147,174.5,-147</points>
<connection>
<GID>197</GID>
<name>N_in0</name></connection>
<intersection>172.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-146.5,172.5,-146.5</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<intersection>172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>220.5,-187,220.5,-156.5</points>
<intersection>-187 1</intersection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210.5,-187,220.5,-187</points>
<connection>
<GID>226</GID>
<name>N_in1</name></connection>
<intersection>220.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220.5,-156.5,230.5,-156.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-165.5,219.5,-154.5</points>
<intersection>-165.5 1</intersection>
<intersection>-154.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-165.5,219.5,-165.5</points>
<connection>
<GID>207</GID>
<name>N_in1</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>219.5,-154.5,230.5,-154.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-152.5,219.5,-142.5</points>
<intersection>-152.5 2</intersection>
<intersection>-142.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,-142.5,219.5,-142.5</points>
<connection>
<GID>192</GID>
<name>N_in1</name></connection>
<intersection>219.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>219.5,-152.5,230.5,-152.5</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>223,-150.5,223,-119.5</points>
<intersection>-150.5 2</intersection>
<intersection>-119.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208.5,-119.5,223,-119.5</points>
<connection>
<GID>243</GID>
<name>N_in1</name></connection>
<intersection>223 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223,-150.5,230.5,-150.5</points>
<connection>
<GID>175</GID>
<name>IN_3</name></connection>
<intersection>223 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>236.5,-153.5,250,-153.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>246</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>169.5,-124,174,-124</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<connection>
<GID>181</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-140,171,-119</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>196</GID>
<name>N_in3</name></connection>
<connection>
<GID>180</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-141.5,193.5,-141.5</points>
<connection>
<GID>188</GID>
<name>N_in1</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>190,-151.5,194,-151.5</points>
<connection>
<GID>189</GID>
<name>N_in1</name></connection>
<connection>
<GID>187</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>200,-150.5,200.5,-150.5</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201.5,-149.5,201.5,-146</points>
<connection>
<GID>190</GID>
<name>N_in3</name></connection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-146,201.5,-146</points>
<intersection>193.5 2</intersection>
<intersection>201.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>193.5,-146,193.5,-143.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>-146 1</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>199.5,-142.5,201,-142.5</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<connection>
<GID>191</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-149.5,191.5,-145</points>
<intersection>-149.5 1</intersection>
<intersection>-145 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-149.5,194,-149.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191.5,-145,202,-145</points>
<intersection>191.5 0</intersection>
<intersection>202 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>202,-145,202,-143.5</points>
<connection>
<GID>191</GID>
<name>N_in2</name></connection>
<intersection>-145 2</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>203,-142.5,207,-142.5</points>
<connection>
<GID>191</GID>
<name>N_in1</name></connection>
<connection>
<GID>192</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>175.5,-153,176,-153</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-141,176,-141</points>
<connection>
<GID>196</GID>
<name>N_in1</name></connection>
<connection>
<GID>193</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-163,171,-142</points>
<connection>
<GID>214</GID>
<name>N_in3</name></connection>
<connection>
<GID>196</GID>
<name>N_in2</name></connection>
<intersection>-153 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>171,-153,171.5,-153</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-146,175.5,-143</points>
<connection>
<GID>197</GID>
<name>N_in3</name></connection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-143,176,-143</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-151,175.5,-148</points>
<connection>
<GID>197</GID>
<name>N_in2</name></connection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-151,176,-151</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-142,185,-141.5</points>
<intersection>-142 2</intersection>
<intersection>-141.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-141.5,188,-141.5</points>
<connection>
<GID>188</GID>
<name>N_in0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182,-142,185,-142</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-152,185,-151.5</points>
<intersection>-152 2</intersection>
<intersection>-151.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-151.5,188,-151.5</points>
<connection>
<GID>189</GID>
<name>N_in0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>182,-152,185,-152</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,-164.5,193,-164.5</points>
<connection>
<GID>203</GID>
<name>N_in1</name></connection>
<connection>
<GID>201</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,-174.5,193.5,-174.5</points>
<connection>
<GID>204</GID>
<name>N_in1</name></connection>
<connection>
<GID>202</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>199.5,-173.5,200,-173.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<connection>
<GID>205</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-172.5,201,-169</points>
<connection>
<GID>205</GID>
<name>N_in3</name></connection>
<intersection>-169 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-169,201,-169</points>
<intersection>193 2</intersection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>193,-169,193,-166.5</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>-169 1</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>199,-165.5,200.5,-165.5</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<connection>
<GID>206</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-172.5,191,-168</points>
<intersection>-172.5 1</intersection>
<intersection>-168 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-172.5,193.5,-172.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-168,201.5,-168</points>
<intersection>191 0</intersection>
<intersection>201.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201.5,-168,201.5,-166.5</points>
<connection>
<GID>206</GID>
<name>N_in2</name></connection>
<intersection>-168 2</intersection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>202.5,-165.5,206.5,-165.5</points>
<connection>
<GID>206</GID>
<name>N_in1</name></connection>
<connection>
<GID>207</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>175,-177,175.5,-177</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>175 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>175,-177,175,-176</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>-177 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-164,175.5,-164</points>
<connection>
<GID>214</GID>
<name>N_in1</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-169,175,-166</points>
<connection>
<GID>215</GID>
<name>N_in3</name></connection>
<intersection>-166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-166,175.5,-166</points>
<connection>
<GID>210</GID>
<name>IN_1</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-175,175,-171</points>
<connection>
<GID>215</GID>
<name>N_in2</name></connection>
<intersection>-175 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-175,175.5,-175</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-165,184.5,-164.5</points>
<intersection>-165 2</intersection>
<intersection>-164.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-164.5,187.5,-164.5</points>
<connection>
<GID>203</GID>
<name>N_in0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-165,184.5,-165</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184.5,-176,184.5,-174.5</points>
<intersection>-176 2</intersection>
<intersection>-174.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184.5,-174.5,187.5,-174.5</points>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<intersection>184.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181.5,-176,184.5,-176</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-186,195,-186</points>
<connection>
<GID>222</GID>
<name>N_in1</name></connection>
<connection>
<GID>220</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>191.5,-196,195.5,-196</points>
<connection>
<GID>223</GID>
<name>N_in1</name></connection>
<connection>
<GID>221</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>201.5,-195,202,-195</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>224</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>203,-198.5,203,-194</points>
<connection>
<GID>224</GID>
<name>N_in3</name></connection>
<intersection>-198.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194,-198.5,203,-198.5</points>
<intersection>194 2</intersection>
<intersection>203 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>194,-198.5,194,-188</points>
<intersection>-198.5 1</intersection>
<intersection>-188 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>194,-188,195,-188</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>194 2</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>201,-187,202.5,-187</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<connection>
<GID>225</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-196,192,-194</points>
<intersection>-196 2</intersection>
<intersection>-194 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-194,195.5,-194</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>192,-196,205,-196</points>
<intersection>192 0</intersection>
<intersection>205 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>205,-196,205,-188</points>
<intersection>-196 2</intersection>
<intersection>-188 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>203.5,-188,205,-188</points>
<connection>
<GID>225</GID>
<name>N_in2</name></connection>
<intersection>205 3</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>204.5,-187,208.5,-187</points>
<connection>
<GID>225</GID>
<name>N_in1</name></connection>
<connection>
<GID>226</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>177,-197.5,177.5,-197.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172,-185.5,177.5,-185.5</points>
<connection>
<GID>231</GID>
<name>N_in1</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-197.5,171.5,-186.5</points>
<intersection>-197.5 8</intersection>
<intersection>-186.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>171,-186.5,171.5,-186.5</points>
<connection>
<GID>231</GID>
<name>N_in2</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>171.5,-197.5,173,-197.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-190.5,177,-187.5</points>
<connection>
<GID>232</GID>
<name>N_in3</name></connection>
<intersection>-187.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-187.5,177.5,-187.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-195.5,177,-192.5</points>
<connection>
<GID>232</GID>
<name>N_in2</name></connection>
<intersection>-195.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-195.5,177.5,-195.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-186.5,186.5,-186</points>
<intersection>-186.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,-186,189.5,-186</points>
<connection>
<GID>222</GID>
<name>N_in0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-186.5,186.5,-186.5</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-196.5,186.5,-196</points>
<intersection>-196.5 2</intersection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186.5,-196,189.5,-196</points>
<connection>
<GID>223</GID>
<name>N_in0</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-196.5,186.5,-196.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,-118.5,193,-118.5</points>
<connection>
<GID>238</GID>
<name>N_in1</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>189.5,-128.5,193.5,-128.5</points>
<connection>
<GID>240</GID>
<name>N_in1</name></connection>
<connection>
<GID>237</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>199.5,-127.5,200,-127.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<connection>
<GID>241</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-126.5,201,-123</points>
<connection>
<GID>241</GID>
<name>N_in3</name></connection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-123,201,-123</points>
<intersection>193 2</intersection>
<intersection>201 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>193,-123,193,-120.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>199,-119.5,200.5,-119.5</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<connection>
<GID>242</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-126.5,191,-122</points>
<intersection>-126.5 1</intersection>
<intersection>-122 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-126.5,193.5,-126.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-122,201.5,-122</points>
<intersection>191 0</intersection>
<intersection>201.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>201.5,-122,201.5,-120.5</points>
<connection>
<GID>242</GID>
<name>N_in2</name></connection>
<intersection>-122 2</intersection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>202.5,-119.5,206.5,-119.5</points>
<connection>
<GID>242</GID>
<name>N_in1</name></connection>
<connection>
<GID>243</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>175,-130,175.5,-130</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>172,-118,175.5,-118</points>
<connection>
<GID>180</GID>
<name>N_in1</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-6.15,-49.8817,47.775,-83.1183</PageViewport>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>18.5,-64.5</position>
<gparam>LABEL_TEXT Can change clock cyle by sliding bar at top (next to play button)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>BB_CLOCK</type>
<position>-3,-54.5</position>
<output>
<ID>CLK</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>272</ID>
<type>GA_LED</type>
<position>7,-54.5</position>
<input>
<ID>N_in0</ID>215 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>BB_CLOCK</type>
<position>23,-68.5</position>
<output>
<ID>CLK</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>284</ID>
<type>GA_LED</type>
<position>46.5,-78.5</position>
<input>
<ID>N_in0</ID>232 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>AA_AND2</type>
<position>32.5,-78.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_TOGGLE</type>
<position>13,-79.5</position>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>17.5,-61</position>
<gparam>LABEL_TEXT Clock and clocked circuits</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,-54.5,6,-54.5</points>
<connection>
<GID>269</GID>
<name>CLK</name></connection>
<connection>
<GID>272</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-78.5,45.5,-78.5</points>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<connection>
<GID>284</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-77.5,28,-68.5</points>
<intersection>-77.5 1</intersection>
<intersection>-68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-77.5,29.5,-77.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-68.5,28,-68.5</points>
<connection>
<GID>282</GID>
<name>CLK</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-79.5,29.5,-79.5</points>
<connection>
<GID>286</GID>
<name>OUT_0</name></connection>
<connection>
<GID>285</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>126.45,11.7875,179.275,-20.771</PageViewport>
<gate>
<ID>387</ID>
<type>AA_LABEL</type>
<position>154.5,1</position>
<gparam>LABEL_TEXT When clock is low (0) output does not change even if  D changes</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>147.5,-9.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>389</ID>
<type>AA_LABEL</type>
<position>161,-3</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>AA_LABEL</type>
<position>163,-15.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>AA_LABEL</type>
<position>154.5,7</position>
<gparam>LABEL_TEXT D Latch with Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>BA_NAND2</type>
<position>166,-5.5</position>
<input>
<ID>IN_0</ID>350 </input>
<input>
<ID>IN_1</ID>353 </input>
<output>
<ID>OUT</ID>354 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>393</ID>
<type>BA_NAND2</type>
<position>166.5,-13.5</position>
<input>
<ID>IN_0</ID>355 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>394</ID>
<type>HA_JUNC_2</type>
<position>158.5,-4.5</position>
<input>
<ID>N_in0</ID>363 </input>
<input>
<ID>N_in1</ID>350 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>395</ID>
<type>HA_JUNC_2</type>
<position>158.5,-14.5</position>
<input>
<ID>N_in0</ID>364 </input>
<input>
<ID>N_in1</ID>351 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>396</ID>
<type>HE_JUNC_4</type>
<position>171,-13.5</position>
<input>
<ID>N_in0</ID>352 </input>
<input>
<ID>N_in3</ID>353 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>HE_JUNC_4</type>
<position>171.5,-5.5</position>
<input>
<ID>N_in0</ID>354 </input>
<input>
<ID>N_in1</ID>356 </input>
<input>
<ID>N_in2</ID>355 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>398</ID>
<type>AA_TOGGLE</type>
<position>139,-4</position>
<output>
<ID>OUT_0</ID>359 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>399</ID>
<type>GA_LED</type>
<position>177.5,-5.5</position>
<input>
<ID>N_in0</ID>356 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_LABEL</type>
<position>136.5,-4</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>BA_NAND2</type>
<position>150.5,-4.5</position>
<input>
<ID>IN_0</ID>358 </input>
<input>
<ID>IN_1</ID>361 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>BA_NAND2</type>
<position>151,-14.5</position>
<input>
<ID>IN_0</ID>362 </input>
<input>
<ID>IN_1</ID>357 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>403</ID>
<type>AE_SMALL_INVERTER</type>
<position>146,-15.5</position>
<input>
<ID>IN_0</ID>360 </input>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>404</ID>
<type>HE_JUNC_4</type>
<position>143,-4</position>
<input>
<ID>N_in0</ID>359 </input>
<input>
<ID>N_in1</ID>358 </input>
<input>
<ID>N_in2</ID>360 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>405</ID>
<type>HE_JUNC_4</type>
<position>145.5,-9.5</position>
<input>
<ID>N_in0</ID>365 </input>
<input>
<ID>N_in2</ID>362 </input>
<input>
<ID>N_in3</ID>361 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>406</ID>
<type>BB_CLOCK</type>
<position>138,-9</position>
<output>
<ID>CLK</ID>365 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_LABEL</type>
<position>134.5,-12</position>
<gparam>LABEL_TEXT Connect Clock to WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>385</ID>
<type>AA_LABEL</type>
<position>152,4</position>
<gparam>LABEL_TEXT Q gets updated only when clock is high (1)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-4.5,163,-4.5</points>
<connection>
<GID>394</GID>
<name>N_in1</name></connection>
<connection>
<GID>392</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>159.5,-14.5,163.5,-14.5</points>
<connection>
<GID>395</GID>
<name>N_in1</name></connection>
<connection>
<GID>393</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>169.5,-13.5,170,-13.5</points>
<connection>
<GID>393</GID>
<name>OUT</name></connection>
<connection>
<GID>396</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-12.5,171,-9</points>
<connection>
<GID>396</GID>
<name>N_in3</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-9,171,-9</points>
<intersection>163 2</intersection>
<intersection>171 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>163,-9,163,-6.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>169,-5.5,170.5,-5.5</points>
<connection>
<GID>392</GID>
<name>OUT</name></connection>
<connection>
<GID>397</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-12.5,161,-8</points>
<intersection>-12.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-12.5,163.5,-12.5</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>161,-8,171.5,-8</points>
<intersection>161 0</intersection>
<intersection>171.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>171.5,-8,171.5,-6.5</points>
<connection>
<GID>397</GID>
<name>N_in2</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>172.5,-5.5,176.5,-5.5</points>
<connection>
<GID>397</GID>
<name>N_in1</name></connection>
<connection>
<GID>399</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>148,-15.5,148,-15.5</points>
<connection>
<GID>402</GID>
<name>IN_1</name></connection>
<connection>
<GID>403</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>144,-3.5,147.5,-3.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>144 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>144,-4,144,-3.5</points>
<connection>
<GID>404</GID>
<name>N_in1</name></connection>
<intersection>-3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>141,-4,142,-4</points>
<connection>
<GID>398</GID>
<name>OUT_0</name></connection>
<connection>
<GID>404</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-15.5,143,-5</points>
<connection>
<GID>404</GID>
<name>N_in2</name></connection>
<intersection>-15.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>143,-15.5,144,-15.5</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-8.5,145.5,-5.5</points>
<connection>
<GID>405</GID>
<name>N_in3</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-5.5,147.5,-5.5</points>
<connection>
<GID>401</GID>
<name>IN_1</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-13.5,145.5,-10.5</points>
<connection>
<GID>405</GID>
<name>N_in2</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-13.5,148,-13.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>153.5,-4.5,157.5,-4.5</points>
<connection>
<GID>394</GID>
<name>N_in0</name></connection>
<connection>
<GID>401</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>154,-14.5,157.5,-14.5</points>
<connection>
<GID>395</GID>
<name>N_in0</name></connection>
<connection>
<GID>402</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-9,144.5,-9</points>
<connection>
<GID>406</GID>
<name>CLK</name></connection>
<intersection>144.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>144.5,-9.5,144.5,-9</points>
<connection>
<GID>405</GID>
<name>N_in0</name></connection>
<intersection>-9 1</intersection></vsegment></shape></wire></page 6>
<page 7>
<PageViewport>678.25,-178.609,770.35,-235.375</PageViewport>
<gate>
<ID>336</ID>
<type>AA_LABEL</type>
<position>708,-194.5</position>
<gparam>LABEL_TEXT Latch 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>AA_LABEL</type>
<position>758.5,-196</position>
<gparam>LABEL_TEXT Latch 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>339</ID>
<type>AA_LABEL</type>
<position>701,-205.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>AA_LABEL</type>
<position>682.5,-195.5</position>
<gparam>LABEL_TEXT Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>343</ID>
<type>BA_NAND2</type>
<position>719,-201.5</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_1</ID>276 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>BA_NAND2</type>
<position>719.5,-209.5</position>
<input>
<ID>IN_0</ID>278 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>HA_JUNC_2</type>
<position>711.5,-200.5</position>
<input>
<ID>N_in0</ID>284 </input>
<input>
<ID>N_in1</ID>273 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>HA_JUNC_2</type>
<position>711.5,-210.5</position>
<input>
<ID>N_in0</ID>285 </input>
<input>
<ID>N_in1</ID>274 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>HE_JUNC_4</type>
<position>724,-209.5</position>
<input>
<ID>N_in0</ID>275 </input>
<input>
<ID>N_in3</ID>276 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>HE_JUNC_4</type>
<position>724.5,-201.5</position>
<input>
<ID>N_in0</ID>277 </input>
<input>
<ID>N_in1</ID>348 </input>
<input>
<ID>N_in2</ID>278 </input>
<input>
<ID>N_in3</ID>349 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AA_TOGGLE</type>
<position>684,-199.5</position>
<output>
<ID>OUT_0</ID>281 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_LABEL</type>
<position>689.5,-195.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>351</ID>
<type>BA_NAND2</type>
<position>701.5,-201</position>
<input>
<ID>IN_0</ID>280 </input>
<input>
<ID>IN_1</ID>283 </input>
<output>
<ID>OUT</ID>284 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>BA_NAND2</type>
<position>701.5,-211</position>
<input>
<ID>IN_0</ID>346 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>285 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_SMALL_INVERTER</type>
<position>692,-212</position>
<input>
<ID>IN_0</ID>282 </input>
<output>
<ID>OUT_0</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>354</ID>
<type>HE_JUNC_4</type>
<position>690,-199.5</position>
<input>
<ID>N_in0</ID>281 </input>
<input>
<ID>N_in1</ID>280 </input>
<input>
<ID>N_in2</ID>282 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>HE_JUNC_4</type>
<position>698,-206</position>
<input>
<ID>N_in2</ID>346 </input>
<input>
<ID>N_in3</ID>283 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>746.5,-207</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>359</ID>
<type>BA_NAND2</type>
<position>760,-203.5</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>BA_NAND2</type>
<position>760,-211.5</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>HA_JUNC_2</type>
<position>753,-202.5</position>
<input>
<ID>N_in0</ID>308 </input>
<input>
<ID>N_in1</ID>286 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>HA_JUNC_2</type>
<position>751,-212.5</position>
<input>
<ID>N_in0</ID>345 </input>
<input>
<ID>N_in1</ID>287 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>HE_JUNC_4</type>
<position>765,-211.5</position>
<input>
<ID>N_in0</ID>288 </input>
<input>
<ID>N_in3</ID>289 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>HE_JUNC_4</type>
<position>764.5,-203.5</position>
<input>
<ID>N_in0</ID>293 </input>
<input>
<ID>N_in1</ID>295 </input>
<input>
<ID>N_in2</ID>294 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>GA_LED</type>
<position>767,-203.5</position>
<input>
<ID>N_in0</ID>295 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_LABEL</type>
<position>738.5,-198.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>367</ID>
<type>BA_NAND2</type>
<position>743,-202.5</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>299 </input>
<output>
<ID>OUT</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>BA_NAND2</type>
<position>744,-212.5</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>369</ID>
<type>AE_SMALL_INVERTER</type>
<position>737.5,-213.5</position>
<input>
<ID>IN_0</ID>298 </input>
<output>
<ID>OUT_0</ID>296 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>370</ID>
<type>HE_JUNC_4</type>
<position>734.5,-201.5</position>
<input>
<ID>N_in0</ID>348 </input>
<input>
<ID>N_in1</ID>297 </input>
<input>
<ID>N_in2</ID>298 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>HE_JUNC_4</type>
<position>739.5,-207</position>
<input>
<ID>N_in0</ID>347 </input>
<input>
<ID>N_in2</ID>307 </input>
<input>
<ID>N_in3</ID>299 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>AE_SMALL_INVERTER</type>
<position>714.5,-219.5</position>
<input>
<ID>IN_0</ID>347 </input>
<output>
<ID>OUT_0</ID>346 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>373</ID>
<type>BB_CLOCK</type>
<position>717,-224.5</position>
<output>
<ID>CLK</ID>347 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>374</ID>
<type>GA_LED</type>
<position>724.5,-196.5</position>
<input>
<ID>N_in2</ID>349 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>375</ID>
<type>AA_LABEL</type>
<position>731,-194</position>
<gparam>LABEL_TEXT Q_intermediate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>376</ID>
<type>AA_LABEL</type>
<position>769,-200.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>AA_LABEL</type>
<position>718.5,-188</position>
<gparam>LABEL_TEXT D Flip-Flop: 2 D Latches</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>712.5,-200.5,716,-200.5</points>
<connection>
<GID>345</GID>
<name>N_in1</name></connection>
<connection>
<GID>343</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>712.5,-210.5,716.5,-210.5</points>
<connection>
<GID>346</GID>
<name>N_in1</name></connection>
<connection>
<GID>344</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>722.5,-209.5,723,-209.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<connection>
<GID>347</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>724,-208.5,724,-205</points>
<connection>
<GID>347</GID>
<name>N_in3</name></connection>
<intersection>-205 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>716,-205,724,-205</points>
<intersection>716 2</intersection>
<intersection>724 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>716,-205,716,-202.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>-205 1</intersection></vsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>722,-201.5,723.5,-201.5</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>348</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>714,-208.5,714,-204</points>
<intersection>-208.5 1</intersection>
<intersection>-204 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>714,-208.5,716.5,-208.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>714 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>714,-204,724.5,-204</points>
<intersection>714 0</intersection>
<intersection>724.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>724.5,-204,724.5,-202.5</points>
<connection>
<GID>348</GID>
<name>N_in2</name></connection>
<intersection>-204 2</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>694,-212,698.5,-212</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<connection>
<GID>352</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>691,-199.5,698.5,-199.5</points>
<connection>
<GID>354</GID>
<name>N_in1</name></connection>
<intersection>698.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>698.5,-200,698.5,-199.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-199.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>686,-199.5,689,-199.5</points>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection>
<connection>
<GID>354</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>690,-212,690,-200.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>354</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,-205,698,-202</points>
<connection>
<GID>355</GID>
<name>N_in3</name></connection>
<intersection>-202 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>698,-202,698.5,-202</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>698 0</intersection></hsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>707.5,-201,707.5,-200.5</points>
<intersection>-201 2</intersection>
<intersection>-200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>707.5,-200.5,710.5,-200.5</points>
<connection>
<GID>345</GID>
<name>N_in0</name></connection>
<intersection>707.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>704.5,-201,707.5,-201</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>707.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>707.5,-211,707.5,-210.5</points>
<intersection>-211 2</intersection>
<intersection>-210.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>707.5,-210.5,710.5,-210.5</points>
<connection>
<GID>346</GID>
<name>N_in0</name></connection>
<intersection>707.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>704.5,-211,707.5,-211</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>707.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>754,-202.5,757,-202.5</points>
<connection>
<GID>361</GID>
<name>N_in1</name></connection>
<connection>
<GID>359</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>752,-212.5,757,-212.5</points>
<connection>
<GID>362</GID>
<name>N_in1</name></connection>
<connection>
<GID>360</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>763,-211.5,764,-211.5</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<connection>
<GID>363</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>765,-210.5,765,-208.5</points>
<connection>
<GID>363</GID>
<name>N_in3</name></connection>
<intersection>-208.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>757,-208.5,765,-208.5</points>
<intersection>757 2</intersection>
<intersection>765 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>757,-208.5,757,-204.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>-208.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>763,-203.5,763.5,-203.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<connection>
<GID>364</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>753.5,-210.5,753.5,-206.5</points>
<intersection>-210.5 1</intersection>
<intersection>-206.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>753.5,-210.5,757,-210.5</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>753.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>753.5,-206.5,764.5,-206.5</points>
<intersection>753.5 0</intersection>
<intersection>764.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>764.5,-206.5,764.5,-204.5</points>
<connection>
<GID>364</GID>
<name>N_in2</name></connection>
<intersection>-206.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>765.5,-203.5,766,-203.5</points>
<connection>
<GID>364</GID>
<name>N_in1</name></connection>
<connection>
<GID>365</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>739.5,-213.5,741,-213.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>735.5,-201.5,740,-201.5</points>
<connection>
<GID>370</GID>
<name>N_in1</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>734.5,-213.5,734.5,-202.5</points>
<connection>
<GID>370</GID>
<name>N_in2</name></connection>
<intersection>-213.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>734.5,-213.5,735.5,-213.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>734.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>739.5,-206,739.5,-203.5</points>
<connection>
<GID>371</GID>
<name>N_in3</name></connection>
<intersection>-203.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>739.5,-203.5,740,-203.5</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>739.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>739.5,-211.5,739.5,-208</points>
<connection>
<GID>371</GID>
<name>N_in2</name></connection>
<intersection>-211.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>739.5,-211.5,741,-211.5</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>739.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>746,-202.5,752,-202.5</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<connection>
<GID>361</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>747,-212.5,750,-212.5</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<connection>
<GID>362</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>698,-219.5,698,-207</points>
<connection>
<GID>355</GID>
<name>N_in2</name></connection>
<intersection>-219.5 2</intersection>
<intersection>-210 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>698,-219.5,712.5,-219.5</points>
<connection>
<GID>372</GID>
<name>OUT_0</name></connection>
<intersection>698 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>698,-210,698.5,-210</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>698 0</intersection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>716.5,-219.5,730.5,-219.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>721.5 9</intersection>
<intersection>730.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>730.5,-219.5,730.5,-207</points>
<intersection>-219.5 1</intersection>
<intersection>-207 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>730.5,-207,738.5,-207</points>
<connection>
<GID>371</GID>
<name>N_in0</name></connection>
<intersection>730.5 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>721.5,-224.5,721.5,-219.5</points>
<intersection>-224.5 12</intersection>
<intersection>-219.5 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>721,-224.5,721.5,-224.5</points>
<connection>
<GID>373</GID>
<name>CLK</name></connection>
<intersection>721.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>725.5,-201.5,733.5,-201.5</points>
<connection>
<GID>348</GID>
<name>N_in1</name></connection>
<connection>
<GID>370</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>724.5,-200.5,724.5,-197.5</points>
<connection>
<GID>348</GID>
<name>N_in3</name></connection>
<connection>
<GID>374</GID>
<name>N_in2</name></connection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>127.65,-95.7552,175.55,-125.278</PageViewport>
<gate>
<ID>408</ID>
<type>AE_DFF_LOW_NT</type>
<position>157,-112.5</position>
<input>
<ID>IN_0</ID>367 </input>
<output>
<ID>OUTINV_0</ID>369 </output>
<output>
<ID>OUT_0</ID>368 </output>
<input>
<ID>clock</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_LABEL</type>
<position>150,-102</position>
<gparam>LABEL_TEXT D Flip Flop Schematic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>AA_TOGGLE</type>
<position>141,-110.5</position>
<output>
<ID>OUT_0</ID>367 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>411</ID>
<type>BB_CLOCK</type>
<position>141.5,-115.5</position>
<output>
<ID>CLK</ID>366 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>412</ID>
<type>GA_LED</type>
<position>174,-110.5</position>
<input>
<ID>N_in0</ID>368 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>AA_LABEL</type>
<position>133.5,-110</position>
<gparam>LABEL_TEXT Input D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>414</ID>
<type>AA_LABEL</type>
<position>148.5,-118</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>AA_LABEL</type>
<position>167.5,-107.5</position>
<gparam>LABEL_TEXT Output Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>416</ID>
<type>AA_LABEL</type>
<position>168,-116</position>
<gparam>LABEL_TEXT Output Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>417</ID>
<type>GA_LED</type>
<position>167,-113.5</position>
<input>
<ID>N_in0</ID>369 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-115.5,145.5,-113.5</points>
<connection>
<GID>411</GID>
<name>CLK</name></connection>
<intersection>-113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145.5,-113.5,154,-113.5</points>
<connection>
<GID>408</GID>
<name>clock</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>143,-110.5,154,-110.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<connection>
<GID>410</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160,-110.5,173,-110.5</points>
<connection>
<GID>408</GID>
<name>OUT_0</name></connection>
<connection>
<GID>412</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>160,-113.5,166,-113.5</points>
<connection>
<GID>408</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>417</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>503.156,-110.825,580.844,-158.708</PageViewport>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>535,-122.5</position>
<gparam>LABEL_TEXT D Flip-flop with write enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AF_DFF_LOW</type>
<position>536,-130.5</position>
<input>
<ID>IN_0</ID>379 </input>
<output>
<ID>OUT_0</ID>378 </output>
<input>
<ID>clock</ID>381 </input>
<input>
<ID>clock_enable</ID>380 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>438</ID>
<type>AA_TOGGLE</type>
<position>527,-127</position>
<output>
<ID>OUT_0</ID>379 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>439</ID>
<type>AA_TOGGLE</type>
<position>526,-133.5</position>
<output>
<ID>OUT_0</ID>380 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>440</ID>
<type>GA_LED</type>
<position>544.5,-128.5</position>
<input>
<ID>N_in0</ID>378 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>BB_CLOCK</type>
<position>518,-130.5</position>
<output>
<ID>CLK</ID>381 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>442</ID>
<type>AA_LABEL</type>
<position>522.5,-126.5</position>
<gparam>LABEL_TEXT Input D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>443</ID>
<type>AA_LABEL</type>
<position>523,-135.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>444</ID>
<type>AA_LABEL</type>
<position>550,-128.5</position>
<gparam>LABEL_TEXT Output Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>378</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>539,-128.5,543.5,-128.5</points>
<connection>
<GID>437</GID>
<name>OUT_0</name></connection>
<connection>
<GID>440</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>531,-128.5,531,-127</points>
<intersection>-128.5 1</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>531,-128.5,533,-128.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>531 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>529,-127,531,-127</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<intersection>531 0</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>530.5,-133.5,530.5,-132.5</points>
<intersection>-133.5 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>530.5,-132.5,533,-132.5</points>
<connection>
<GID>437</GID>
<name>clock_enable</name></connection>
<intersection>530.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>528,-133.5,530.5,-133.5</points>
<connection>
<GID>439</GID>
<name>OUT_0</name></connection>
<intersection>530.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>522,-130.5,533,-130.5</points>
<connection>
<GID>441</GID>
<name>CLK</name></connection>
<connection>
<GID>437</GID>
<name>clock</name></connection></hsegment></shape></wire></page 9></circuit>