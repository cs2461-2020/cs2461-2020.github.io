<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>22.8077,-219.475,174.142,-312.75</PageViewport>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>118,-310.5</position>
<gparam>LABEL_TEXT 4-1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>66,-282.5</position>
<gparam>LABEL_TEXT Input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_REGISTER4</type>
<position>99.5,-268</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>52 </output>
<output>
<ID>OUT_1</ID>45 </output>
<output>
<ID>OUT_2</ID>41 </output>
<output>
<ID>OUT_3</ID>37 </output>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>62 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_REGISTER4</type>
<position>99.5,-280.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>51 </output>
<output>
<ID>OUT_1</ID>46 </output>
<output>
<ID>OUT_2</ID>42 </output>
<output>
<ID>OUT_3</ID>38 </output>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>63 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_REGISTER4</type>
<position>99.5,-292.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>50 </output>
<output>
<ID>OUT_1</ID>47 </output>
<output>
<ID>OUT_2</ID>43 </output>
<output>
<ID>OUT_3</ID>39 </output>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>64 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_REGISTER4</type>
<position>99.5,-304.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>57 </input>
<output>
<ID>OUT_0</ID>49 </output>
<output>
<ID>OUT_1</ID>48 </output>
<output>
<ID>OUT_2</ID>44 </output>
<output>
<ID>OUT_3</ID>40 </output>
<input>
<ID>clock</ID>61 </input>
<input>
<ID>load</ID>65 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_MUX_4x1</type>
<position>116.5,-302.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<input>
<ID>SEL_0</ID>67 </input>
<input>
<ID>SEL_1</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>30</ID>
<type>DD_KEYPAD_HEX</type>
<position>80,-240.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<output>
<ID>OUT_1</ID>69 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_MUX_4x1</type>
<position>139,-257</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<output>
<ID>OUT</ID>73 </output>
<input>
<ID>SEL_0</ID>70 </input>
<input>
<ID>SEL_1</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_MUX_4x1</type>
<position>139,-268</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>45 </input>
<output>
<ID>OUT</ID>72 </output>
<input>
<ID>SEL_0</ID>70 </input>
<input>
<ID>SEL_1</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_MUX_4x1</type>
<position>139,-279.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>52 </input>
<output>
<ID>OUT</ID>71 </output>
<input>
<ID>SEL_0</ID>70 </input>
<input>
<ID>SEL_1</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_MUX_4x1</type>
<position>139,-245.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>74 </output>
<input>
<ID>SEL_0</ID>70 </input>
<input>
<ID>SEL_1</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>35</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>151,-265.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>68,-234</position>
<gparam>LABEL_TEXT Address 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>90.5,-220.5</position>
<gparam>LABEL_TEXT What is this circuit? What does it do ?</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AE_MUX_4x1</type>
<position>116.5,-292</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<input>
<ID>IN_2</ID>46 </input>
<input>
<ID>IN_3</ID>45 </input>
<output>
<ID>OUT</ID>54 </output>
<input>
<ID>SEL_0</ID>67 </input>
<input>
<ID>SEL_1</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_MUX_4x1</type>
<position>116,-279.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>41 </input>
<output>
<ID>OUT</ID>55 </output>
<input>
<ID>SEL_0</ID>67 </input>
<input>
<ID>SEL_1</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>40</ID>
<type>AE_MUX_4x1</type>
<position>116,-268.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>38 </input>
<input>
<ID>IN_3</ID>37 </input>
<output>
<ID>OUT</ID>56 </output>
<input>
<ID>SEL_0</ID>67 </input>
<input>
<ID>SEL_1</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>41</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>147.5,-290</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>56 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 6</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>42</ID>
<type>DD_KEYPAD_HEX</type>
<position>76.5,-283</position>
<output>
<ID>OUT_0</ID>60 </output>
<output>
<ID>OUT_1</ID>59 </output>
<output>
<ID>OUT_2</ID>58 </output>
<output>
<ID>OUT_3</ID>57 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>43</ID>
<type>BB_CLOCK</type>
<position>79.5,-310.5</position>
<output>
<ID>CLK</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>61.5,-258</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>BA_DECODER_2x4</type>
<position>85,-259</position>
<input>
<ID>ENABLE</ID>68 </input>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT_0</ID>65 </output>
<output>
<ID>OUT_1</ID>64 </output>
<output>
<ID>OUT_2</ID>63 </output>
<output>
<ID>OUT_3</ID>62 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>DD_KEYPAD_HEX</type>
<position>65.5,-250</position>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>66 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>51.5,-247.5</position>
<gparam>LABEL_TEXT Address 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>54,-260.5</position>
<gparam>LABEL_TEXT Write Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>81,-263</position>
<gparam>LABEL_TEXT 2-4 Decoder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-266,106,-265.5</points>
<intersection>-266 2</intersection>
<intersection>-265.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-265.5,127.5,-265.5</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<intersection>106 0</intersection>
<intersection>127.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-266,106,-266</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>106 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>127.5,-265.5,127.5,-242.5</points>
<intersection>-265.5 1</intersection>
<intersection>-242.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>127.5,-242.5,136,-242.5</points>
<connection>
<GID>34</GID>
<name>IN_3</name></connection>
<intersection>127.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-278.5,106,-267.5</points>
<intersection>-278.5 2</intersection>
<intersection>-267.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-267.5,128,-267.5</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<intersection>106 0</intersection>
<intersection>128 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-278.5,106,-278.5</points>
<connection>
<GID>26</GID>
<name>OUT_3</name></connection>
<intersection>106 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-267.5,128,-244.5</points>
<intersection>-267.5 1</intersection>
<intersection>-244.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128,-244.5,136,-244.5</points>
<connection>
<GID>34</GID>
<name>IN_2</name></connection>
<intersection>128 3</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-290.5,106.5,-269.5</points>
<intersection>-290.5 2</intersection>
<intersection>-269.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-269.5,128,-269.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>106.5 0</intersection>
<intersection>128 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-290.5,106.5,-290.5</points>
<connection>
<GID>27</GID>
<name>OUT_3</name></connection>
<intersection>106.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128,-269.5,128,-246.5</points>
<intersection>-269.5 1</intersection>
<intersection>-246.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128,-246.5,136,-246.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>128 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-302.5,107,-271.5</points>
<intersection>-302.5 2</intersection>
<intersection>-271.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-271.5,128.5,-271.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection>
<intersection>128.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-302.5,107,-302.5</points>
<connection>
<GID>28</GID>
<name>OUT_3</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-271.5,128.5,-248.5</points>
<intersection>-271.5 1</intersection>
<intersection>-248.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128.5,-248.5,136,-248.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>128.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-276.5,129,-254</points>
<intersection>-276.5 1</intersection>
<intersection>-254 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-276.5,129,-276.5</points>
<connection>
<GID>39</GID>
<name>IN_3</name></connection>
<intersection>103.5 4</intersection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129,-254,136,-254</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>129 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>103.5,-276.5,103.5,-267</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>-276.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-279.5,107.5,-278.5</points>
<intersection>-279.5 2</intersection>
<intersection>-278.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-278.5,130,-278.5</points>
<connection>
<GID>39</GID>
<name>IN_2</name></connection>
<intersection>107.5 0</intersection>
<intersection>130 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-279.5,107.5,-279.5</points>
<connection>
<GID>26</GID>
<name>OUT_2</name></connection>
<intersection>107.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>130,-278.5,130,-256</points>
<intersection>-278.5 1</intersection>
<intersection>-256 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>130,-256,136,-256</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>130 3</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-291.5,107.5,-280.5</points>
<intersection>-291.5 2</intersection>
<intersection>-280.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-280.5,130.5,-280.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>107.5 0</intersection>
<intersection>130.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-291.5,107.5,-291.5</points>
<connection>
<GID>27</GID>
<name>OUT_2</name></connection>
<intersection>107.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>130.5,-280.5,130.5,-258</points>
<intersection>-280.5 1</intersection>
<intersection>-258 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>130.5,-258,136,-258</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>130.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-303.5,108,-282.5</points>
<intersection>-303.5 1</intersection>
<intersection>-282.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-303.5,108,-303.5</points>
<connection>
<GID>28</GID>
<name>OUT_2</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108,-282.5,131,-282.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection>
<intersection>131 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131,-282.5,131,-260</points>
<intersection>-282.5 2</intersection>
<intersection>-260 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>131,-260,136,-260</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>131 3</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-289,109,-268</points>
<intersection>-289 2</intersection>
<intersection>-268 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-268,109,-268</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>109 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>109,-289,131.5,-289</points>
<connection>
<GID>38</GID>
<name>IN_3</name></connection>
<intersection>109 0</intersection>
<intersection>131.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>131.5,-289,131.5,-265</points>
<intersection>-289 2</intersection>
<intersection>-265 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>131.5,-265,136,-265</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<intersection>131.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-291,109.5,-281</points>
<intersection>-291 1</intersection>
<intersection>-281 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-291,132,-291</points>
<connection>
<GID>38</GID>
<name>IN_2</name></connection>
<intersection>109.5 0</intersection>
<intersection>132 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-281,109.5,-281</points>
<intersection>103.5 3</intersection>
<intersection>109.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103.5,-281,103.5,-280.5</points>
<connection>
<GID>26</GID>
<name>OUT_1</name></connection>
<intersection>-281 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>132,-291,132,-267</points>
<intersection>-291 1</intersection>
<intersection>-267 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>132,-267,136,-267</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>132 6</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-293,108.5,-292.5</points>
<intersection>-293 1</intersection>
<intersection>-292.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-293,132.5,-293</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>108.5 0</intersection>
<intersection>132.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-292.5,108.5,-292.5</points>
<connection>
<GID>27</GID>
<name>OUT_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132.5,-293,132.5,-269</points>
<intersection>-293 1</intersection>
<intersection>-269 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>132.5,-269,136,-269</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>132.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-304.5,108.5,-295</points>
<intersection>-304.5 2</intersection>
<intersection>-295 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-295,133,-295</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection>
<intersection>133 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-304.5,108.5,-304.5</points>
<connection>
<GID>28</GID>
<name>OUT_1</name></connection>
<intersection>108.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133,-295,133,-271</points>
<intersection>-295 1</intersection>
<intersection>-271 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>133,-271,136,-271</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>133 3</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-305.5,136,-305.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>136 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>136,-305.5,136,-282.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-305.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-304.5,110,-296.5</points>
<intersection>-304.5 5</intersection>
<intersection>-303.5 2</intersection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-296.5,110,-296.5</points>
<intersection>103.5 3</intersection>
<intersection>110 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-303.5,113.5,-303.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>110 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103.5,-296.5,103.5,-293.5</points>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection>
<intersection>-296.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>110,-304.5,135.5,-304.5</points>
<intersection>110 0</intersection>
<intersection>135.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>135.5,-304.5,135.5,-280.5</points>
<intersection>-304.5 5</intersection>
<intersection>-280.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>135.5,-280.5,136,-280.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>135.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-301.5,111,-281.5</points>
<intersection>-301.5 4</intersection>
<intersection>-281.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>103.5,-281.5,111,-281.5</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>111 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>111,-301.5,135,-301.5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>111 0</intersection>
<intersection>135 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>135,-301.5,135,-278.5</points>
<intersection>-301.5 4</intersection>
<intersection>-278.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>135,-278.5,136,-278.5</points>
<connection>
<GID>33</GID>
<name>IN_2</name></connection>
<intersection>135 6</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-299.5,112,-269</points>
<intersection>-299.5 2</intersection>
<intersection>-269 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-269,112,-269</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>112,-299.5,134.5,-299.5</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<intersection>112 0</intersection>
<intersection>134.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>134.5,-299.5,134.5,-276.5</points>
<intersection>-299.5 2</intersection>
<intersection>-276.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>134.5,-276.5,136,-276.5</points>
<connection>
<GID>33</GID>
<name>IN_3</name></connection>
<intersection>134.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-302.5,125,-291</points>
<intersection>-302.5 1</intersection>
<intersection>-291 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119.5,-302.5,125,-302.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,-291,144.5,-291</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-292,123.5,-290</points>
<intersection>-292 2</intersection>
<intersection>-290 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-290,144.5,-290</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-292,123.5,-292</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-289,123.5,-279.5</points>
<intersection>-289 2</intersection>
<intersection>-279.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-279.5,123.5,-279.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-289,144.5,-289</points>
<connection>
<GID>41</GID>
<name>IN_2</name></connection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-288,124.5,-268.5</points>
<intersection>-288 2</intersection>
<intersection>-268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>119,-268.5,124.5,-268.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-288,144.5,-288</points>
<connection>
<GID>41</GID>
<name>IN_3</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-280,81.5,-266</points>
<connection>
<GID>42</GID>
<name>OUT_3</name></connection>
<intersection>-278.5 3</intersection>
<intersection>-266 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-266,95.5,-266</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81.5,-278.5,95.5,-278.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>81.5 0</intersection>
<intersection>93 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93,-302.5,93,-278.5</points>
<intersection>-302.5 7</intersection>
<intersection>-290.5 5</intersection>
<intersection>-278.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>93,-290.5,95.5,-290.5</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>93 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>93,-302.5,95.5,-302.5</points>
<connection>
<GID>28</GID>
<name>IN_3</name></connection>
<intersection>93 4</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-282,84.5,-267</points>
<intersection>-282 2</intersection>
<intersection>-279.5 3</intersection>
<intersection>-267 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-267,95.5,-267</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-282,84.5,-282</points>
<connection>
<GID>42</GID>
<name>OUT_2</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>84.5,-279.5,95.5,-279.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>84.5 0</intersection>
<intersection>94 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>94,-303.5,94,-279.5</points>
<intersection>-303.5 7</intersection>
<intersection>-291.5 5</intersection>
<intersection>-279.5 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>94,-291.5,95.5,-291.5</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>94 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>94,-303.5,95.5,-303.5</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>94 4</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-292.5,88.5,-268</points>
<intersection>-292.5 4</intersection>
<intersection>-284 2</intersection>
<intersection>-280.5 3</intersection>
<intersection>-268 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88.5,-268,95.5,-268</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-284,88.5,-284</points>
<connection>
<GID>42</GID>
<name>OUT_1</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-280.5,95.5,-280.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>88.5,-292.5,95.5,-292.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>88.5 0</intersection>
<intersection>92 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>92,-304.5,92,-292.5</points>
<intersection>-304.5 6</intersection>
<intersection>-292.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>92,-304.5,95.5,-304.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>92 5</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-305.5,90.5,-269</points>
<intersection>-305.5 6</intersection>
<intersection>-293.5 4</intersection>
<intersection>-286 2</intersection>
<intersection>-281.5 3</intersection>
<intersection>-269 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-269,95.5,-269</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-286,90.5,-286</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>90.5,-281.5,95.5,-281.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>90.5,-293.5,95.5,-293.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>90.5,-305.5,95.5,-305.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-310.5,85,-296.5</points>
<intersection>-310.5 1</intersection>
<intersection>-308.5 4</intersection>
<intersection>-296.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-310.5,85,-310.5</points>
<connection>
<GID>43</GID>
<name>CLK</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>85,-296.5,98.5,-296.5</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>85 0</intersection>
<intersection>85.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>85,-308.5,98.5,-308.5</points>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>85.5,-296.5,85.5,-272</points>
<intersection>-296.5 3</intersection>
<intersection>-284.5 6</intersection>
<intersection>-272 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>85.5,-284.5,98.5,-284.5</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>85.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>85.5,-272,98.5,-272</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>85.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-263,98.5,-257.5</points>
<connection>
<GID>25</GID>
<name>load</name></connection>
<intersection>-257.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-257.5,98.5,-257.5</points>
<connection>
<GID>45</GID>
<name>OUT_3</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-275.5,95,-258.5</points>
<intersection>-275.5 2</intersection>
<intersection>-258.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-258.5,95,-258.5</points>
<connection>
<GID>45</GID>
<name>OUT_2</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95,-275.5,98.5,-275.5</points>
<connection>
<GID>26</GID>
<name>load</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-287.5,94.5,-259.5</points>
<intersection>-287.5 2</intersection>
<intersection>-259.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-259.5,94.5,-259.5</points>
<connection>
<GID>45</GID>
<name>OUT_1</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-287.5,98.5,-287.5</points>
<connection>
<GID>27</GID>
<name>load</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-299.5,96,-260.5</points>
<intersection>-299.5 2</intersection>
<intersection>-260.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-260.5,96,-260.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96,-299.5,98.5,-299.5</points>
<connection>
<GID>28</GID>
<name>load</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-251,121.5,-251</points>
<connection>
<GID>46</GID>
<name>OUT_1</name></connection>
<intersection>71.5 6</intersection>
<intersection>121.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>121.5,-296.5,121.5,-251</points>
<intersection>-296.5 18</intersection>
<intersection>-287 19</intersection>
<intersection>-273.5 14</intersection>
<intersection>-262.5 10</intersection>
<intersection>-251 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>71.5,-259.5,71.5,-251</points>
<intersection>-259.5 7</intersection>
<intersection>-251 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>71.5,-259.5,82,-259.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>71.5 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>116,-262.5,121.5,-262.5</points>
<intersection>116 12</intersection>
<intersection>121.5 5</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>116,-274.5,116,-262.5</points>
<connection>
<GID>39</GID>
<name>SEL_1</name></connection>
<connection>
<GID>40</GID>
<name>SEL_1</name></connection>
<intersection>-273.5 14</intersection>
<intersection>-262.5 10</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>116,-273.5,121.5,-273.5</points>
<intersection>116 12</intersection>
<intersection>121.5 5</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>116.5,-296.5,121.5,-296.5</points>
<intersection>116.5 20</intersection>
<intersection>121.5 5</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>116.5,-287,121.5,-287</points>
<connection>
<GID>38</GID>
<name>SEL_1</name></connection>
<intersection>121.5 5</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>116.5,-297.5,116.5,-296.5</points>
<connection>
<GID>29</GID>
<name>SEL_1</name></connection>
<intersection>-296.5 18</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-260.5,70.5,-253</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>-260.5 5</intersection>
<intersection>-253 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-253,119.5,-253</points>
<intersection>70.5 0</intersection>
<intersection>119.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>119.5,-297.5,119.5,-253</points>
<intersection>-297.5 12</intersection>
<intersection>-287 10</intersection>
<intersection>-274.5 7</intersection>
<intersection>-263.5 8</intersection>
<intersection>-253 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>70.5,-260.5,82,-260.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>117,-274.5,119.5,-274.5</points>
<connection>
<GID>39</GID>
<name>SEL_0</name></connection>
<intersection>119.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>117,-263.5,119.5,-263.5</points>
<connection>
<GID>40</GID>
<name>SEL_0</name></connection>
<intersection>119.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>117.5,-287,119.5,-287</points>
<connection>
<GID>38</GID>
<name>SEL_0</name></connection>
<intersection>119.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>117.5,-297.5,119.5,-297.5</points>
<connection>
<GID>29</GID>
<name>SEL_0</name></connection>
<intersection>119.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-257.5,82,-257.5</points>
<connection>
<GID>45</GID>
<name>ENABLE</name></connection>
<intersection>64.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64.5,-258,64.5,-257.5</points>
<intersection>-258 4</intersection>
<intersection>-257.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-258,64.5,-258</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>64.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-274.5,139,-240.5</points>
<connection>
<GID>34</GID>
<name>SEL_1</name></connection>
<connection>
<GID>33</GID>
<name>SEL_1</name></connection>
<connection>
<GID>32</GID>
<name>SEL_1</name></connection>
<connection>
<GID>31</GID>
<name>SEL_1</name></connection>
<intersection>-247.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-247.5,139,-247.5</points>
<intersection>87 12</intersection>
<intersection>139 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>87,-247.5,87,-241.5</points>
<intersection>-247.5 1</intersection>
<intersection>-241.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>85,-241.5,87,-241.5</points>
<connection>
<GID>30</GID>
<name>OUT_1</name></connection>
<intersection>87 12</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-274.5,140,-240.5</points>
<connection>
<GID>34</GID>
<name>SEL_0</name></connection>
<connection>
<GID>33</GID>
<name>SEL_0</name></connection>
<connection>
<GID>32</GID>
<name>SEL_0</name></connection>
<connection>
<GID>31</GID>
<name>SEL_0</name></connection>
<intersection>-249.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-249.5,140,-249.5</points>
<intersection>87 2</intersection>
<intersection>140 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>87,-249.5,87,-243.5</points>
<intersection>-249.5 1</intersection>
<intersection>-243.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>85,-243.5,87,-243.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>87 2</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-279.5,145,-266.5</points>
<intersection>-279.5 2</intersection>
<intersection>-266.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-266.5,148,-266.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-279.5,145,-279.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>142,-265.5,148,-265.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>142 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>142,-268,142,-265.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>-265.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-264.5,145,-257</points>
<intersection>-264.5 2</intersection>
<intersection>-257 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-257,145,-257</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,-264.5,148,-264.5</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-263.5,146.5,-245.5</points>
<intersection>-263.5 2</intersection>
<intersection>-245.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-245.5,146.5,-245.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-263.5,148,-263.5</points>
<connection>
<GID>35</GID>
<name>IN_3</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>328.942,265.525,559.858,123.2</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>392.5,264.5</position>
<gparam>LABEL_TEXT What is this circuit? What does it do ?</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_REGISTER4</type>
<position>424.5,189.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT_0</ID>10 </output>
<output>
<ID>OUT_1</ID>11 </output>
<output>
<ID>OUT_2</ID>12 </output>
<output>
<ID>OUT_3</ID>13 </output>
<input>
<ID>clock</ID>9 </input>
<input>
<ID>load</ID>35 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_REGISTER4</type>
<position>424.5,167.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT_0</ID>17 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>15 </output>
<output>
<ID>OUT_3</ID>14 </output>
<input>
<ID>clock</ID>9 </input>
<input>
<ID>load</ID>36 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>4</ID>
<type>DD_KEYPAD_HEX</type>
<position>398.5,189.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<output>
<ID>OUT_1</ID>3 </output>
<output>
<ID>OUT_2</ID>2 </output>
<output>
<ID>OUT_3</ID>1 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>5</ID>
<type>DD_KEYPAD_HEX</type>
<position>397.5,167.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<output>
<ID>OUT_1</ID>7 </output>
<output>
<ID>OUT_2</ID>6 </output>
<output>
<ID>OUT_3</ID>5 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BB_CLOCK</type>
<position>412.5,136.5</position>
<output>
<ID>CLK</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_FULLADDER_4BIT</type>
<position>463.5,178.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>14 </input>
<input>
<ID>IN_B_0</ID>10 </input>
<input>
<ID>IN_B_1</ID>11 </input>
<input>
<ID>IN_B_2</ID>12 </input>
<input>
<ID>IN_B_3</ID>13 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>26 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>28 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>8</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>465,141.5</position>
<output>
<ID>A_equal_B</ID>23 </output>
<output>
<ID>A_greater_B</ID>22 </output>
<output>
<ID>A_less_B</ID>24 </output>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>14 </input>
<input>
<ID>IN_B_0</ID>10 </input>
<input>
<ID>IN_B_1</ID>11 </input>
<input>
<ID>IN_B_2</ID>12 </input>
<input>
<ID>IN_B_3</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>426,184.5</position>
<gparam>LABEL_TEXT Number Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>428,162</position>
<gparam>LABEL_TEXT Number X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>461.5,189.5</position>
<gparam>LABEL_TEXT Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>439,125</position>
<gparam>LABEL_TEXT Compare: out=4 if Y>X, 1 if X >Y, 0 if X=Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_MUX_2x1</type>
<position>482,175</position>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>21 </output>
<input>
<ID>SEL_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_MUX_2x1</type>
<position>482,166</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>20 </output>
<input>
<ID>SEL_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_MUX_2x1</type>
<position>482,157</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>19 </output>
<input>
<ID>SEL_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_MUX_2x1</type>
<position>482,147.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>18 </output>
<input>
<ID>SEL_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>504.5,160.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>20 </input>
<input>
<ID>IN_3</ID>21 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_ROM_4x4</type>
<position>383,244.5</position>
<input>
<ID>ADDRESS_0</ID>33 </input>
<input>
<ID>ADDRESS_1</ID>32 </input>
<input>
<ID>ADDRESS_2</ID>31 </input>
<input>
<ID>ADDRESS_3</ID>30 </input>
<output>
<ID>DATA_OUT_0</ID>35 </output>
<output>
<ID>DATA_OUT_1</ID>36 </output>
<output>
<ID>DATA_OUT_2</ID>29 </output>
<input>
<ID>ENABLE_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 4</lparam></gate>
<gate>
<ID>19</ID>
<type>DD_KEYPAD_HEX</type>
<position>358.5,244</position>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>30 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>400,244</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>355.5,251.5</position>
<gparam>LABEL_TEXT Address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>407.5,238.5</position>
<gparam>LABEL_TEXT Output - contents at address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>433.5,259</position>
<gparam>LABEL_TEXT The "program" in memory determines which function is 'called'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>451,255</position>
<gparam>LABEL_TEXT The output of ROM sets the control lines: determines which register is written into and which function implemented</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,191.5,412,192.5</points>
<intersection>191.5 1</intersection>
<intersection>192.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>412,191.5,420.5,191.5</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403.5,192.5,412,192.5</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>403.5,190.5,420.5,190.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,188.5,412,189.5</points>
<intersection>188.5 1</intersection>
<intersection>189.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403.5,188.5,412,188.5</points>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,189.5,420.5,189.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>412,186.5,412,188.5</points>
<intersection>186.5 1</intersection>
<intersection>188.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>403.5,186.5,412,186.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>412 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>412,188.5,420.5,188.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>412 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411.5,169.5,411.5,170.5</points>
<intersection>169.5 1</intersection>
<intersection>170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>411.5,169.5,420.5,169.5</points>
<connection>
<GID>3</GID>
<name>IN_3</name></connection>
<intersection>411.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>402.5,170.5,411.5,170.5</points>
<connection>
<GID>5</GID>
<name>OUT_3</name></connection>
<intersection>411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>402.5,168.5,420.5,168.5</points>
<connection>
<GID>5</GID>
<name>OUT_2</name></connection>
<connection>
<GID>3</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411.5,166.5,411.5,167.5</points>
<intersection>166.5 1</intersection>
<intersection>167.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,166.5,411.5,166.5</points>
<connection>
<GID>5</GID>
<name>OUT_1</name></connection>
<intersection>411.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>411.5,167.5,420.5,167.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>411.5,164.5,411.5,166.5</points>
<intersection>164.5 1</intersection>
<intersection>166.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,164.5,411.5,164.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>411.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>411.5,166.5,420.5,166.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>418.5,136.5,418.5,185.5</points>
<intersection>136.5 1</intersection>
<intersection>163.5 3</intersection>
<intersection>185.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>416.5,136.5,418.5,136.5</points>
<connection>
<GID>6</GID>
<name>CLK</name></connection>
<intersection>418.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>418.5,185.5,423.5,185.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>418.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>418.5,163.5,423.5,163.5</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>418.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,183.5,444,188.5</points>
<intersection>183.5 2</intersection>
<intersection>188.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,188.5,444,188.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,183.5,461,183.5</points>
<connection>
<GID>7</GID>
<name>IN_B_0</name></connection>
<intersection>444 0</intersection>
<intersection>461 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>461,146.5,461,183.5</points>
<connection>
<GID>8</GID>
<name>IN_B_0</name></connection>
<intersection>183.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445.5,182.5,445.5,189.5</points>
<intersection>182.5 2</intersection>
<intersection>189.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,189.5,445.5,189.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>445.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>445.5,182.5,461,182.5</points>
<connection>
<GID>7</GID>
<name>IN_B_1</name></connection>
<intersection>445.5 0</intersection>
<intersection>461 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>461,145.5,461,182.5</points>
<connection>
<GID>8</GID>
<name>IN_B_1</name></connection>
<intersection>182.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>446.5,181.5,446.5,190.5</points>
<intersection>181.5 2</intersection>
<intersection>190.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,190.5,446.5,190.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>446.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>446.5,181.5,461,181.5</points>
<connection>
<GID>7</GID>
<name>IN_B_2</name></connection>
<intersection>446.5 0</intersection>
<intersection>461 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>461,144.5,461,181.5</points>
<connection>
<GID>8</GID>
<name>IN_B_2</name></connection>
<intersection>181.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445,180.5,445,191.5</points>
<intersection>180.5 2</intersection>
<intersection>191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,191.5,445,191.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>445 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>445,180.5,461,180.5</points>
<connection>
<GID>7</GID>
<name>IN_B_3</name></connection>
<intersection>445 0</intersection>
<intersection>461 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>461,143.5,461,180.5</points>
<connection>
<GID>8</GID>
<name>IN_B_3</name></connection>
<intersection>180.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,169.5,444,173.5</points>
<intersection>169.5 1</intersection>
<intersection>173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,169.5,444,169.5</points>
<connection>
<GID>3</GID>
<name>OUT_3</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,173.5,461,173.5</points>
<connection>
<GID>7</GID>
<name>IN_3</name></connection>
<intersection>444 0</intersection>
<intersection>461 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>461,136.5,461,173.5</points>
<connection>
<GID>8</GID>
<name>IN_3</name></connection>
<intersection>173.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>445,137.5,445,174.5</points>
<intersection>137.5 3</intersection>
<intersection>168.5 1</intersection>
<intersection>174.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,168.5,445,168.5</points>
<connection>
<GID>3</GID>
<name>OUT_2</name></connection>
<intersection>445 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>445,174.5,459.5,174.5</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>445 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>445,137.5,461,137.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>445 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444,138.5,444,175.5</points>
<intersection>138.5 3</intersection>
<intersection>167.5 1</intersection>
<intersection>175.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,167.5,444,167.5</points>
<connection>
<GID>3</GID>
<name>OUT_1</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444,175.5,459.5,175.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>444 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>444,138.5,461,138.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>444 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>446,139.5,446,176.5</points>
<intersection>139.5 3</intersection>
<intersection>166.5 1</intersection>
<intersection>176.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,166.5,446,166.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>446 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>446,176.5,459.5,176.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>446 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>446,139.5,461,139.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>446 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,147.5,492.5,159.5</points>
<intersection>147.5 1</intersection>
<intersection>159.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,147.5,492.5,147.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,159.5,501.5,159.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,157,492.5,160.5</points>
<intersection>157 1</intersection>
<intersection>160.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,157,492.5,157</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,160.5,501.5,160.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,161.5,492.5,166</points>
<intersection>161.5 2</intersection>
<intersection>166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,166,492.5,166</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,161.5,501.5,161.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>492.5,162.5,492.5,175</points>
<intersection>162.5 2</intersection>
<intersection>175 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>484,175,492.5,175</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>492.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>492.5,162.5,501.5,162.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>492.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,128,463,133.5</points>
<connection>
<GID>8</GID>
<name>A_greater_B</name></connection>
<intersection>128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>463,128,480,128</points>
<intersection>463 0</intersection>
<intersection>480 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>480,128,480,146.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>128 1</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>465,129,465,133.5</points>
<connection>
<GID>8</GID>
<name>A_equal_B</name></connection>
<intersection>129 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>465,129,477.5,129</points>
<intersection>465 0</intersection>
<intersection>477.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>477.5,129,477.5,156</points>
<intersection>129 1</intersection>
<intersection>156 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>477.5,156,480,156</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>477.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>475.5,133.5,475.5,165</points>
<intersection>133.5 2</intersection>
<intersection>165 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>475.5,165,480,165</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>475.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>467,133.5,475.5,133.5</points>
<connection>
<GID>8</GID>
<name>A_less_B</name></connection>
<intersection>475.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>471,148.5,471,180</points>
<intersection>148.5 2</intersection>
<intersection>180 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,180,471,180</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>471 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>471,148.5,480,148.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>471 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,158,469.5,179</points>
<intersection>158 2</intersection>
<intersection>179 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,179,469.5,179</points>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection>
<intersection>469.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>469.5,158,480,158</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>469.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>472,167,472,178</points>
<intersection>167 2</intersection>
<intersection>178 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,178,472,178</points>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection>
<intersection>472 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>472,167,480,167</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>472 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>473.5,176,473.5,177</points>
<intersection>176 2</intersection>
<intersection>177 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>467.5,177,473.5,177</points>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection>
<intersection>473.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>473.5,176,480,176</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>473.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>487.5,150,487.5,230.5</points>
<intersection>150 4</intersection>
<intersection>159.5 5</intersection>
<intersection>168.5 6</intersection>
<intersection>177.5 7</intersection>
<intersection>230.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>382.5,230.5,487.5,230.5</points>
<intersection>382.5 3</intersection>
<intersection>487.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>382.5,230.5,382.5,239.5</points>
<connection>
<GID>18</GID>
<name>DATA_OUT_2</name></connection>
<intersection>230.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>482,150,487.5,150</points>
<connection>
<GID>16</GID>
<name>SEL_0</name></connection>
<intersection>487.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>482,159.5,487.5,159.5</points>
<connection>
<GID>15</GID>
<name>SEL_0</name></connection>
<intersection>487.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>482,168.5,487.5,168.5</points>
<connection>
<GID>14</GID>
<name>SEL_0</name></connection>
<intersection>487.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>482,177.5,487.5,177.5</points>
<connection>
<GID>13</GID>
<name>SEL_0</name></connection>
<intersection>487.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>364,246,364,247</points>
<intersection>246 3</intersection>
<intersection>247 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>364,246,378,246</points>
<connection>
<GID>18</GID>
<name>ADDRESS_3</name></connection>
<intersection>364 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>363.5,247,364,247</points>
<connection>
<GID>19</GID>
<name>OUT_3</name></connection>
<intersection>364 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>363.5,245,378,245</points>
<connection>
<GID>18</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>19</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365.5,243,365.5,244</points>
<intersection>243 2</intersection>
<intersection>244 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>363.5,243,365.5,243</points>
<connection>
<GID>19</GID>
<name>OUT_1</name></connection>
<intersection>365.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>365.5,244,378,244</points>
<connection>
<GID>18</GID>
<name>ADDRESS_1</name></connection>
<intersection>365.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>366.5,241,366.5,243</points>
<intersection>241 2</intersection>
<intersection>243 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>363.5,241,366.5,241</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>366.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>366.5,243,378,243</points>
<connection>
<GID>18</GID>
<name>ADDRESS_0</name></connection>
<intersection>366.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>388,244,398,244</points>
<connection>
<GID>18</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,217,384.5,239.5</points>
<connection>
<GID>18</GID>
<name>DATA_OUT_0</name></connection>
<intersection>217 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>423.5,194.5,423.5,217</points>
<connection>
<GID>2</GID>
<name>load</name></connection>
<intersection>217 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>384.5,217,423.5,217</points>
<intersection>384.5 0</intersection>
<intersection>423.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>383.5,206,383.5,239.5</points>
<connection>
<GID>18</GID>
<name>DATA_OUT_1</name></connection>
<intersection>206 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>414.5,172.5,414.5,206</points>
<intersection>172.5 3</intersection>
<intersection>206 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>383.5,206,414.5,206</points>
<intersection>383.5 0</intersection>
<intersection>414.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>414.5,172.5,423.5,172.5</points>
<connection>
<GID>3</GID>
<name>load</name></connection>
<intersection>414.5 1</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-125.55,37.7665,87.1001,-93.3</PageViewport>
<gate>
<ID>50</ID>
<type>AA_REGISTER4</type>
<position>-11.5,-27</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>77 </input>
<input>
<ID>IN_2</ID>76 </input>
<input>
<ID>IN_3</ID>75 </input>
<output>
<ID>OUT_0</ID>84 </output>
<output>
<ID>OUT_1</ID>85 </output>
<output>
<ID>OUT_2</ID>86 </output>
<output>
<ID>OUT_3</ID>87 </output>
<input>
<ID>clock</ID>83 </input>
<input>
<ID>load</ID>105 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_REGISTER4</type>
<position>-11.5,-49</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>80 </input>
<input>
<ID>IN_3</ID>79 </input>
<output>
<ID>OUT_0</ID>91 </output>
<output>
<ID>OUT_1</ID>90 </output>
<output>
<ID>OUT_2</ID>89 </output>
<output>
<ID>OUT_3</ID>88 </output>
<input>
<ID>clock</ID>83 </input>
<input>
<ID>load</ID>106 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>52</ID>
<type>DD_KEYPAD_HEX</type>
<position>-37.5,-26.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<output>
<ID>OUT_1</ID>77 </output>
<output>
<ID>OUT_2</ID>76 </output>
<output>
<ID>OUT_3</ID>75 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>53</ID>
<type>DD_KEYPAD_HEX</type>
<position>-38.5,-49</position>
<output>
<ID>OUT_0</ID>82 </output>
<output>
<ID>OUT_1</ID>81 </output>
<output>
<ID>OUT_2</ID>80 </output>
<output>
<ID>OUT_3</ID>79 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>54</ID>
<type>BB_CLOCK</type>
<position>-23.5,-80</position>
<output>
<ID>CLK</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_FULLADDER_4BIT</type>
<position>27.5,-38</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>88 </input>
<input>
<ID>IN_B_0</ID>84 </input>
<input>
<ID>IN_B_1</ID>85 </input>
<input>
<ID>IN_B_2</ID>86 </input>
<input>
<ID>IN_B_3</ID>87 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>100 </output>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_3</ID>102 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>56</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>29,-75</position>
<output>
<ID>A_equal_B</ID>97 </output>
<output>
<ID>A_greater_B</ID>96 </output>
<output>
<ID>A_less_B</ID>98 </output>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>89 </input>
<input>
<ID>IN_3</ID>88 </input>
<input>
<ID>IN_B_0</ID>84 </input>
<input>
<ID>IN_B_1</ID>85 </input>
<input>
<ID>IN_B_2</ID>86 </input>
<input>
<ID>IN_B_3</ID>87 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>-10,-32</position>
<gparam>LABEL_TEXT Number Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>-8,-54.5</position>
<gparam>LABEL_TEXT Number X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>25.5,-27</position>
<gparam>LABEL_TEXT Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>3,-91.5</position>
<gparam>LABEL_TEXT Compare: out=4 if Y>X, 1 if X >Y, 0 if X=Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_MUX_2x1</type>
<position>46,-41.5</position>
<input>
<ID>IN_1</ID>102 </input>
<output>
<ID>OUT</ID>95 </output>
<input>
<ID>SEL_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_MUX_2x1</type>
<position>46,-50.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>94 </output>
<input>
<ID>SEL_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_MUX_2x1</type>
<position>46,-59.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>93 </output>
<input>
<ID>SEL_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_MUX_2x1</type>
<position>46,-69</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>92 </output>
<input>
<ID>SEL_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>68.5,-56</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>93 </input>
<input>
<ID>IN_2</ID>94 </input>
<input>
<ID>IN_3</ID>95 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>66</ID>
<type>BA_ROM_4x4</type>
<position>-53,28</position>
<input>
<ID>ADDRESS_0</ID>108 </input>
<input>
<ID>ADDRESS_1</ID>113 </input>
<input>
<ID>ADDRESS_2</ID>114 </input>
<input>
<ID>ADDRESS_3</ID>115 </input>
<output>
<ID>DATA_OUT_0</ID>105 </output>
<output>
<ID>DATA_OUT_1</ID>106 </output>
<output>
<ID>DATA_OUT_2</ID>103 </output>
<input>
<ID>ENABLE_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:1 1</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:3 4</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>-36,27.5</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>-102,15</position>
<gparam>LABEL_TEXT Address</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-29,18.5</position>
<gparam>LABEL_TEXT Output - contents at address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_REGISTER4</type>
<position>-80,7.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>111 </input>
<input>
<ID>IN_2</ID>112 </input>
<input>
<ID>IN_3</ID>110 </input>
<output>
<ID>OUT_0</ID>108 </output>
<output>
<ID>OUT_1</ID>113 </output>
<output>
<ID>OUT_2</ID>114 </output>
<output>
<ID>OUT_3</ID>115 </output>
<input>
<ID>clock</ID>83 </input>
<input>
<ID>count_enable</ID>107 </input>
<input>
<ID>count_up</ID>107 </input>
<input>
<ID>load</ID>116 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>-93.5,17</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>72</ID>
<type>DD_KEYPAD_HEX</type>
<position>-102,6.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>112 </output>
<output>
<ID>OUT_3</ID>110 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>-71.5,1</position>
<gparam>LABEL_TEXT Register Counts up</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>-100.5,19.5</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>-94,22.5</position>
<gparam>LABEL_TEXT Load initial address</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>-56.5,37</position>
<gparam>LABEL_TEXT Similar to Page2...But address incremented each cycle in ROM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-25,-24,-23.5</points>
<intersection>-25 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-25,-15.5,-25</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>-24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-23.5,-24,-23.5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32.5,-25.5,-15.5,-25.5</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>-15.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-15.5,-26,-15.5,-25.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32.5,-27.5,-15.5,-27.5</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>-15.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15.5,-27.5,-15.5,-27</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-29.5,-24,-28</points>
<intersection>-29.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-32.5,-29.5,-24,-29.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>-24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24,-28,-15.5,-28</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-47,-24.5,-46</points>
<intersection>-47 1</intersection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-47,-15.5,-47</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33.5,-46,-24.5,-46</points>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33.5,-48,-15.5,-48</points>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection>
<connection>
<GID>51</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-50,-24.5,-49</points>
<intersection>-50 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-50,-24.5,-50</points>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-49,-15.5,-49</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-52,-24.5,-50</points>
<intersection>-52 1</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,-52,-24.5,-52</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-50,-15.5,-50</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-80,-17.5,-31</points>
<intersection>-80 1</intersection>
<intersection>-76 6</intersection>
<intersection>-53 3</intersection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-80,-17.5,-80</points>
<connection>
<GID>54</GID>
<name>CLK</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-17.5,-31,-12.5,-31</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17.5,-53,-12.5,-53</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-81,-76,-17.5,-76</points>
<intersection>-81 7</intersection>
<intersection>-17.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-81,-76,-81,3.5</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>-76 6</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-33,8,-28</points>
<intersection>-33 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-28,8,-28</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-33,25,-33</points>
<connection>
<GID>55</GID>
<name>IN_B_0</name></connection>
<intersection>8 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-70,25,-33</points>
<connection>
<GID>56</GID>
<name>IN_B_0</name></connection>
<intersection>-33 2</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-34,8,-27</points>
<intersection>-34 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-27,8,-27</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-34,25,-34</points>
<connection>
<GID>55</GID>
<name>IN_B_1</name></connection>
<intersection>8 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-71,25,-34</points>
<connection>
<GID>56</GID>
<name>IN_B_1</name></connection>
<intersection>-34 2</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-35,8,-26</points>
<intersection>-35 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-26,8,-26</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-35,25,-35</points>
<connection>
<GID>55</GID>
<name>IN_B_2</name></connection>
<intersection>8 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-72,25,-35</points>
<connection>
<GID>56</GID>
<name>IN_B_2</name></connection>
<intersection>-35 2</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-36,8,-25</points>
<intersection>-36 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-25,8,-25</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-36,25,-36</points>
<connection>
<GID>55</GID>
<name>IN_B_3</name></connection>
<intersection>8 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-73,25,-36</points>
<connection>
<GID>56</GID>
<name>IN_B_3</name></connection>
<intersection>-36 2</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-47,8,-43</points>
<intersection>-47 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-47,8,-47</points>
<connection>
<GID>51</GID>
<name>OUT_3</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-43,25,-43</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<intersection>8 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-80,25,-43</points>
<connection>
<GID>56</GID>
<name>IN_3</name></connection>
<intersection>-43 2</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-79,8,-42</points>
<intersection>-79 3</intersection>
<intersection>-48 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-48,8,-48</points>
<connection>
<GID>51</GID>
<name>OUT_2</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-42,23.5,-42</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-79,25,-79</points>
<connection>
<GID>56</GID>
<name>IN_2</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-78,8,-41</points>
<intersection>-78 3</intersection>
<intersection>-49 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-49,8,-49</points>
<connection>
<GID>51</GID>
<name>OUT_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-41,23.5,-41</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-78,25,-78</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-77,8,-40</points>
<intersection>-77 3</intersection>
<intersection>-50 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-50,8,-50</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-40,23.5,-40</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-77,25,-77</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-69,56.5,-57</points>
<intersection>-69 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-69,56.5,-69</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-57,65.5,-57</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-59.5,56.5,-56</points>
<intersection>-59.5 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-59.5,56.5,-59.5</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-56,65.5,-56</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-55,56.5,-50.5</points>
<intersection>-55 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-50.5,56.5,-50.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-55,65.5,-55</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-54,56.5,-41.5</points>
<intersection>-54 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-41.5,56.5,-41.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-54,65.5,-54</points>
<connection>
<GID>65</GID>
<name>IN_3</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-88.5,27,-83</points>
<connection>
<GID>56</GID>
<name>A_greater_B</name></connection>
<intersection>-88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-88.5,44,-88.5</points>
<intersection>27 0</intersection>
<intersection>44 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>44,-88.5,44,-70</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-88.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-87.5,29,-83</points>
<connection>
<GID>56</GID>
<name>A_equal_B</name></connection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-87.5,41.5,-87.5</points>
<intersection>29 0</intersection>
<intersection>41.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>41.5,-87.5,41.5,-60.5</points>
<intersection>-87.5 1</intersection>
<intersection>-60.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>41.5,-60.5,44,-60.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>41.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-83,39.5,-51.5</points>
<intersection>-83 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-51.5,44,-51.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-83,39.5,-83</points>
<connection>
<GID>56</GID>
<name>A_less_B</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-68,37.5,-36.5</points>
<intersection>-68 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-36.5,37.5,-36.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-68,44,-68</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-58.5,37.5,-37.5</points>
<intersection>-58.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-37.5,37.5,-37.5</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-58.5,44,-58.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-49.5,37.5,-38.5</points>
<intersection>-49.5 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-38.5,37.5,-38.5</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-49.5,44,-49.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-40.5,37.5,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-39.5,37.5,-39.5</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-40.5,44,-40.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-66.5,51.5,14</points>
<intersection>-66.5 4</intersection>
<intersection>-57 5</intersection>
<intersection>-48 6</intersection>
<intersection>-39 7</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,14,51.5,14</points>
<intersection>-53.5 3</intersection>
<intersection>51.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-53.5,14,-53.5,23</points>
<connection>
<GID>66</GID>
<name>DATA_OUT_2</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46,-66.5,51.5,-66.5</points>
<connection>
<GID>64</GID>
<name>SEL_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>46,-57,51.5,-57</points>
<connection>
<GID>63</GID>
<name>SEL_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>46,-48,51.5,-48</points>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>46,-39,51.5,-39</points>
<connection>
<GID>61</GID>
<name>SEL_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-48,27.5,-38,27.5</points>
<connection>
<GID>66</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,0.5,-51.5,23</points>
<connection>
<GID>66</GID>
<name>DATA_OUT_0</name></connection>
<intersection>0.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-12.5,-22,-12.5,0.5</points>
<connection>
<GID>50</GID>
<name>load</name></connection>
<intersection>0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-51.5,0.5,-12.5,0.5</points>
<intersection>-51.5 0</intersection>
<intersection>-12.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,-10.5,-52.5,23</points>
<connection>
<GID>66</GID>
<name>DATA_OUT_1</name></connection>
<intersection>-10.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-21.5,-44,-21.5,-10.5</points>
<intersection>-44 3</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-10.5,-21.5,-10.5</points>
<intersection>-52.5 0</intersection>
<intersection>-21.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-21.5,-44,-12.5,-44</points>
<connection>
<GID>51</GID>
<name>load</name></connection>
<intersection>-21.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80,12.5,-80,17</points>
<connection>
<GID>70</GID>
<name>count_enable</name></connection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-91.5,17,-79,17</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-80 0</intersection>
<intersection>-79 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-79,12.5,-79,17</points>
<connection>
<GID>70</GID>
<name>count_up</name></connection>
<intersection>17 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,6.5,-63.5,26.5</points>
<intersection>6.5 2</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,26.5,-58,26.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_0</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,6.5,-63.5,6.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89.5,3.5,-89.5,6.5</points>
<intersection>3.5 2</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-89.5,6.5,-84,6.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,3.5,-89.5,3.5</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,9.5,-84,9.5</points>
<connection>
<GID>72</GID>
<name>OUT_3</name></connection>
<connection>
<GID>70</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90.5,5.5,-90.5,7.5</points>
<intersection>5.5 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-90.5,7.5,-84,7.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,5.5,-90.5,5.5</points>
<connection>
<GID>72</GID>
<name>OUT_1</name></connection>
<intersection>-90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-90.5,7.5,-90.5,8.5</points>
<intersection>7.5 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-90.5,8.5,-84,8.5</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>-90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-97,7.5,-90.5,7.5</points>
<connection>
<GID>72</GID>
<name>OUT_2</name></connection>
<intersection>-90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,7.5,-65,27.5</points>
<intersection>7.5 2</intersection>
<intersection>27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,27.5,-58,27.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_1</name></connection>
<intersection>-65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,7.5,-65,7.5</points>
<connection>
<GID>70</GID>
<name>OUT_1</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66,8.5,-66,28.5</points>
<intersection>8.5 2</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66,28.5,-58,28.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_2</name></connection>
<intersection>-66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,8.5,-66,8.5</points>
<connection>
<GID>70</GID>
<name>OUT_2</name></connection>
<intersection>-66 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,9.5,-67,29.5</points>
<intersection>9.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,29.5,-58,29.5</points>
<connection>
<GID>66</GID>
<name>ADDRESS_3</name></connection>
<intersection>-67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,9.5,-67,9.5</points>
<connection>
<GID>70</GID>
<name>OUT_3</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,12.5,-81,19.5</points>
<connection>
<GID>70</GID>
<name>load</name></connection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98.5,19.5,-81,19.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-81 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>116.835,271.456,1474.83,-565.544</PageViewport></page 3>
<page 4>
<PageViewport>71.9122,400.99,1429.91,-436.01</PageViewport></page 4>
<page 5>
<PageViewport>161.65,664.494,1519.65,-172.506</PageViewport></page 5>
<page 6>
<PageViewport>185.383,700.384,1543.38,-136.616</PageViewport></page 6>
<page 7>
<PageViewport>269.664,436.812,1627.66,-400.188</PageViewport></page 7>
<page 8>
<PageViewport>76.8415,257.28,1434.84,-579.72</PageViewport></page 8>
<page 9>
<PageViewport>591.278,336.427,1949.28,-500.573</PageViewport></page 9></circuit>