<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-35.9,29.683,37.7,-15.6801</PageViewport>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>-2.5,5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>-3,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>-20,6.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>-20,2.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>5,5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>5,-4</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-24.5,6.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>-24,2.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>10.5,5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>9,-4</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>1,19.5</position>
<gparam>LABEL_TEXT What are the truth tables for S0, C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>-9,15</position>
<gparam>LABEL_TEXT What function is this ?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,6,-12,6.5</points>
<intersection>6 1</intersection>
<intersection>6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,6,-5.5,6</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection>
<intersection>-9.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,6.5,-12,6.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-9.5,-3,-9.5,6</points>
<intersection>-3 4</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-9.5,-3,-6,-3</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-9.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-5,-12,4</points>
<intersection>-5 4</intersection>
<intersection>2.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,4,-5.5,4</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,2.5,-12,2.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-12,-5,-6,-5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,5,4,5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<connection>
<GID>11</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-4,4,-4</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>13</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>105.005,4.65776,230.538,-72.7144</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>162,-24</position>
<gparam>LABEL_TEXT C0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>165.5,-6</position>
<gparam>LABEL_TEXT Inputs: A0, B0, C0   Outputs: X0, Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>168,-61</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>144,-11.5</position>
<gparam>LABEL_TEXT What does this circuit do</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AI_XOR2</type>
<position>159,-34.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>141.5,-33</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>141.5,-37</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>137,-33</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>137.5,-37</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>177.5,-33.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>166.5,-26</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>153.5,-46</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>170.5,-46</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>162.5,-54.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>186,-33.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>162.5,-61</position>
<input>
<ID>N_in3</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>192.5,-34</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>162.5,-15</position>
<gparam>LABEL_TEXT Observe how this circuit is built using the circuit from page 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>140,-18</position>
<gparam>LABEL_TEXT (2 Page 1 circuits are combined)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-33.5,149.5,-33</points>
<intersection>-33.5 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-33.5,156,-33.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection>
<intersection>152.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-33,149.5,-33</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>152.5,-43,152.5,-33.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-43,154.5,-35.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-37 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154.5,-35.5,156,-35.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-37,154.5,-37</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162,-34.5,174.5,-34.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>169.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>169.5,-43,169.5,-34.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171.5,-43,171.5,-26</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171.5,-32.5,174.5,-32.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>171.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168.5,-26,171.5,-26</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-50.5,153.5,-49</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>161.5,-51.5,161.5,-50.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>153.5,-50.5,161.5,-50.5</points>
<intersection>153.5 0</intersection>
<intersection>161.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-50.5,170.5,-49</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>163.5,-51.5,163.5,-50.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>163.5,-50.5,170.5,-50.5</points>
<intersection>163.5 1</intersection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>180.5,-33.5,185,-33.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162.5,-60,162.5,-57.5</points>
<connection>
<GID>33</GID>
<name>N_in3</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>184.557,-52.4122,435.643,-207.168</PageViewport>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>265.5,-87.5</position>
<gparam>LABEL_TEXT Observe similarity to Circuit on Page 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>260,-97.5</position>
<gparam>LABEL_TEXT This input C0 is always =0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AI_XOR2</type>
<position>282.5,-110</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>265,-108.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>265,-112.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>260.5,-108.5</position>
<gparam>LABEL_TEXT A0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>261,-112.5</position>
<gparam>LABEL_TEXT B0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AI_XOR2</type>
<position>301,-109</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>290,-101.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>277,-121.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>294,-121.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_OR2</type>
<position>286,-130</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>309.5,-109</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>316,-109.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>291.5,-136.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AI_XOR2</type>
<position>274,-156.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>256.5,-155</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>256.5,-159</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>252,-155</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>252.5,-159</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AI_XOR2</type>
<position>292.5,-155.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND2</type>
<position>268.5,-168</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>285.5,-168</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_OR2</type>
<position>277.5,-176.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>GA_LED</type>
<position>301,-155.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>277.5,-183</position>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>273.5,-147.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>283,-183</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>257,-72.5</position>
<gparam>LABEL_TEXT What is this circuit?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>253.5,-81.5</position>
<gparam>LABEL_TEXT Inputs: A0,A1, B0,B1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>292,-81</position>
<gparam>LABEL_TEXT Outputs:  X0,X1,Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>307.5,-154.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>278.5,-186</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>306.5,-73</position>
<gparam>LABEL_TEXT What "function" is being computed?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>251,-134.5</position>
<gparam>LABEL_TEXT (Page 2 circuit is replicated twice here)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>243.5,-141.5</position>
<gparam>LABEL_TEXT (Output from one Page 2 circuit is input to next one)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>283,-101</position>
<gparam>LABEL_TEXT C0= 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-109,273,-108.5</points>
<intersection>-109 1</intersection>
<intersection>-108.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273,-109,279.5,-109</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection>
<intersection>276 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>267,-108.5,273,-108.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>273 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>276,-118.5,276,-109</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-112.5,273,-111</points>
<intersection>-112.5 2</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273,-111,279.5,-111</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>273 0</intersection>
<intersection>278 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>267,-112.5,273,-112.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>273 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>278,-118.5,278,-111</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-111 1</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>285.5,-110,298,-110</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>293 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>293,-118.5,293,-110</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-110 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-118.5,295,-101.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-108 1</intersection>
<intersection>-101.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295,-108,298,-108</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>292,-101.5,295,-101.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-126,277,-124.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-126 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>285,-127,285,-126</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>277,-126,285,-126</points>
<intersection>277 0</intersection>
<intersection>285 1</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-126,294,-124.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-126 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>287,-127,287,-126</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-126 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>287,-126,294,-126</points>
<intersection>287 1</intersection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>304,-109,308.5,-109</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-155.5,264.5,-155</points>
<intersection>-155.5 1</intersection>
<intersection>-155 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-155.5,271,-155.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>264.5 0</intersection>
<intersection>267.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>258.5,-155,264.5,-155</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>267.5,-165,267.5,-155.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-155.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-159,264.5,-157.5</points>
<intersection>-159 2</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264.5,-157.5,271,-157.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>264.5 0</intersection>
<intersection>269.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>258.5,-159,264.5,-159</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>264.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>269.5,-165,269.5,-157.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268.5,-172.5,268.5,-171</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>-172.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>276.5,-173.5,276.5,-172.5</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>268.5,-172.5,276.5,-172.5</points>
<intersection>268.5 0</intersection>
<intersection>276.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>285.5,-172.5,285.5,-171</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-172.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>278.5,-173.5,278.5,-172.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>278.5,-172.5,285.5,-172.5</points>
<intersection>278.5 1</intersection>
<intersection>285.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>295.5,-155.5,300,-155.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-165,286.5,-149</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-154.5 3</intersection>
<intersection>-149 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>286,-149,286,-133</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>-149 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>286,-149,286.5,-149</points>
<intersection>286 1</intersection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286.5,-154.5,289.5,-154.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277,-156.5,289.5,-156.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>284.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>284.5,-165,284.5,-156.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-156.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-182,277.5,-179.5</points>
<connection>
<GID>59</GID>
<name>N_in3</name></connection>
<connection>
<GID>57</GID>
<name>OUT</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-286.112,85.0057,-49.0885,-61.0829</PageViewport>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-190.5,-30</position>
<gparam>LABEL_TEXT 4-bit input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>-191.5,-25.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>-151.5,-29.5</position>
<gparam>LABEL_TEXT 4-bit input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>-161,21</position>
<input>
<ID>N_in2</ID>46 </input>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>-148,21</position>
<input>
<ID>N_in2</ID>45 </input>
<input>
<ID>N_in3</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>-175.5,66</position>
<gparam>LABEL_TEXT 4-bit Full Adder: Chaining multiple 1-bit adders</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>-174.5,13</position>
<gparam>LABEL_TEXT Output Sum bits</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-149,18</position>
<gparam>LABEL_TEXT bit 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>-206.5,22</position>
<gparam>LABEL_TEXT Overflow?</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-123.5,0.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>48 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 7</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_FULLADDER_1BIT</type>
<position>-148,27</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_B_0</ID>35 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>carry_in</ID>30 </input>
<output>
<ID>carry_out</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_FULLADDER_1BIT</type>
<position>-161,27</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_B_0</ID>36 </input>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>carry_in</ID>29 </input>
<output>
<ID>carry_out</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_FULLADDER_1BIT</type>
<position>-172.5,27</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_B_0</ID>37 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>carry_in</ID>28 </input>
<output>
<ID>carry_out</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_FULLADDER_1BIT</type>
<position>-185.5,27</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_B_0</ID>38 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>carry_in</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>FF_GND</type>
<position>-139.5,26</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>DD_KEYPAD_HEX</type>
<position>-200.5,57.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>33 </output>
<output>
<ID>OUT_3</ID>34 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>80</ID>
<type>DD_KEYPAD_HEX</type>
<position>-201,43.5</position>
<output>
<ID>OUT_0</ID>35 </output>
<output>
<ID>OUT_1</ID>36 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>38 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 5</lparam></gate>
<gate>
<ID>81</ID>
<type>HE_JUNC_4</type>
<position>-179.5,27</position>
<input>
<ID>N_in0</ID>40 </input>
<input>
<ID>N_in1</ID>39 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>-185.5,21</position>
<input>
<ID>N_in0</ID>48 </input>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>-172.5,21</position>
<input>
<ID>N_in2</ID>47 </input>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-167,-38</position>
<gparam>LABEL_TEXT 4-bit output displayed in hex</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-152,-26</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-170.5,-34</position>
<gparam>LABEL_TEXT (X+Y)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>-163,-17</position>
<gparam>LABEL_TEXT Carry-in=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>-148,62.5</position>
<gparam>LABEL_TEXT Carry out from bit i goes to carry-in of bit i+1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>-136,28</position>
<gparam>LABEL_TEXT C0=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>-143,32</position>
<gparam>LABEL_TEXT bit 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>-210.5,59.5</position>
<gparam>LABEL_TEXT Keypad </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-213.5,55.5</position>
<gparam>LABEL_TEXT 4-bit (Hex)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-191.5,31.5</position>
<gparam>LABEL_TEXT bit 3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-175.5,-20</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<input>
<ID>IN_2</ID>128 </input>
<input>
<ID>IN_3</ID>129 </input>
<input>
<ID>IN_B_0</ID>110 </input>
<input>
<ID>IN_B_1</ID>111 </input>
<input>
<ID>IN_B_2</ID>112 </input>
<input>
<ID>IN_B_3</ID>116 </input>
<output>
<ID>OUT_0</ID>130 </output>
<output>
<ID>OUT_1</ID>131 </output>
<output>
<ID>OUT_2</ID>132 </output>
<output>
<ID>OUT_3</ID>133 </output>
<input>
<ID>carry_in</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>-173.5,-8</position>
<gparam>LABEL_TEXT Schematic for 4-bit Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>FF_GND</type>
<position>-164.5,-20.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>147</ID>
<type>DD_KEYPAD_HEX</type>
<position>-191.5,-17.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<output>
<ID>OUT_1</ID>127 </output>
<output>
<ID>OUT_2</ID>128 </output>
<output>
<ID>OUT_3</ID>129 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>153</ID>
<type>DD_KEYPAD_HEX</type>
<position>-153,-18.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_1</ID>111 </output>
<output>
<ID>OUT_2</ID>112 </output>
<output>
<ID>OUT_3</ID>116 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 4</lparam></gate>
<gate>
<ID>184</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-169.5,-28.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>131 </input>
<input>
<ID>IN_2</ID>132 </input>
<input>
<ID>IN_3</ID>133 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 10</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>-191.5,48</position>
<gparam>LABEL_TEXT bit 3 (MSB)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>-192,39.5</position>
<gparam>LABEL_TEXT bit 0 (LSB)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-168.5,27,-165,27</points>
<connection>
<GID>76</GID>
<name>carry_in</name></connection>
<connection>
<GID>75</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,27,-152,27</points>
<connection>
<GID>75</GID>
<name>carry_in</name></connection>
<connection>
<GID>74</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-144,27,-139.5,27</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>74</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-147,30,-147,54.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195.5,54.5,-147,54.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-147 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-160,30,-160,56.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195.5,56.5,-160,56.5</points>
<connection>
<GID>79</GID>
<name>OUT_1</name></connection>
<intersection>-160 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-171.5,30,-171.5,58.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195.5,58.5,-171.5,58.5</points>
<connection>
<GID>79</GID>
<name>OUT_2</name></connection>
<intersection>-171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-184.5,30,-184.5,60.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-195.5,60.5,-184.5,60.5</points>
<connection>
<GID>79</GID>
<name>OUT_3</name></connection>
<intersection>-184.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-149,30,-149,40.5</points>
<connection>
<GID>74</GID>
<name>IN_B_0</name></connection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196,40.5,-149,40.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-149 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-162,30,-162,42.5</points>
<connection>
<GID>75</GID>
<name>IN_B_0</name></connection>
<intersection>42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196,42.5,-162,42.5</points>
<connection>
<GID>80</GID>
<name>OUT_1</name></connection>
<intersection>-162 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-173.5,30,-173.5,44.5</points>
<connection>
<GID>76</GID>
<name>IN_B_0</name></connection>
<intersection>44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196,44.5,-173.5,44.5</points>
<connection>
<GID>80</GID>
<name>OUT_2</name></connection>
<intersection>-173.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-186.5,30,-186.5,46.5</points>
<connection>
<GID>77</GID>
<name>IN_B_0</name></connection>
<intersection>46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196,46.5,-186.5,46.5</points>
<connection>
<GID>80</GID>
<name>OUT_3</name></connection>
<intersection>-186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-178.5,27,-176.5,27</points>
<connection>
<GID>81</GID>
<name>N_in1</name></connection>
<connection>
<GID>76</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-181.5,27,-180.5,27</points>
<connection>
<GID>77</GID>
<name>carry_in</name></connection>
<connection>
<GID>81</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-185.5,22,-185.5,24</points>
<connection>
<GID>82</GID>
<name>N_in3</name></connection>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-172.5,22,-172.5,24</points>
<connection>
<GID>83</GID>
<name>N_in3</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-161,22,-161,24</points>
<connection>
<GID>67</GID>
<name>N_in3</name></connection>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148,22,-148,24</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-148,-0.5,-148,20</points>
<connection>
<GID>68</GID>
<name>N_in2</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-148,-0.5,-126.5,-0.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-148 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-161,0.5,-161,20</points>
<connection>
<GID>67</GID>
<name>N_in2</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-161,0.5,-126.5,0.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-161 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-172.5,1.5,-172.5,20</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-172.5,1.5,-126.5,1.5</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>-172.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-156.5,2.5,-156.5,21</points>
<intersection>2.5 2</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-186.5,21,-156.5,21</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<intersection>-156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-156.5,2.5,-126.5,2.5</points>
<connection>
<GID>73</GID>
<name>IN_3</name></connection>
<intersection>-156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-164.5,-19.5,-164.5,-19</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-167.5,-19,-164.5,-19</points>
<connection>
<GID>131</GID>
<name>carry_in</name></connection>
<intersection>-164.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-170.5,-16,-170.5,-10</points>
<connection>
<GID>131</GID>
<name>IN_B_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-170.5,-10,-143.5,-10</points>
<intersection>-170.5 0</intersection>
<intersection>-143.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-143.5,-21.5,-143.5,-10</points>
<intersection>-21.5 3</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-148,-21.5,-143.5,-21.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>-143.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-171.5,-16,-171.5,-10.5</points>
<connection>
<GID>131</GID>
<name>IN_B_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-171.5,-10.5,-144.5,-10.5</points>
<intersection>-171.5 0</intersection>
<intersection>-144.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-144.5,-19.5,-144.5,-10.5</points>
<intersection>-19.5 3</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-148,-19.5,-144.5,-19.5</points>
<connection>
<GID>153</GID>
<name>OUT_1</name></connection>
<intersection>-144.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-172.5,-16,-172.5,-11</points>
<connection>
<GID>131</GID>
<name>IN_B_2</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-172.5,-11,-146,-11</points>
<intersection>-172.5 0</intersection>
<intersection>-146 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-146,-17.5,-146,-11</points>
<intersection>-17.5 3</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-148,-17.5,-146,-17.5</points>
<connection>
<GID>153</GID>
<name>OUT_2</name></connection>
<intersection>-146 2</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-173.5,-16,-173.5,-11.5</points>
<connection>
<GID>131</GID>
<name>IN_B_3</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-173.5,-11.5,-148,-11.5</points>
<intersection>-173.5 0</intersection>
<intersection>-148 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-148,-15.5,-148,-11.5</points>
<connection>
<GID>153</GID>
<name>OUT_3</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177.5,-16,-177.5,-10</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-184,-10,-177.5,-10</points>
<intersection>-184 2</intersection>
<intersection>-177.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-184,-20.5,-184,-10</points>
<intersection>-20.5 3</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-186.5,-20.5,-184,-20.5</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>-184 2</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178.5,-16,-178.5,-10.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-185,-10.5,-178.5,-10.5</points>
<intersection>-185 2</intersection>
<intersection>-178.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-185,-18.5,-185,-10.5</points>
<intersection>-18.5 3</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-186.5,-18.5,-185,-18.5</points>
<connection>
<GID>147</GID>
<name>OUT_1</name></connection>
<intersection>-185 2</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-179.5,-16,-179.5,-11</points>
<connection>
<GID>131</GID>
<name>IN_2</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-185.5,-11,-179.5,-11</points>
<intersection>-185.5 2</intersection>
<intersection>-179.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-185.5,-16.5,-185.5,-11</points>
<intersection>-16.5 3</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-186.5,-16.5,-185.5,-16.5</points>
<connection>
<GID>147</GID>
<name>OUT_2</name></connection>
<intersection>-185.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-180.5,-16,-180.5,-14.5</points>
<connection>
<GID>131</GID>
<name>IN_3</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-186.5,-14.5,-180.5,-14.5</points>
<connection>
<GID>147</GID>
<name>OUT_3</name></connection>
<intersection>-180.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-174,-29.5,-174,-24</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-174,-29.5,-172.5,-29.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-174 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-175,-28.5,-175,-24</points>
<connection>
<GID>131</GID>
<name>OUT_1</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-175,-28.5,-172.5,-28.5</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>-175 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-176,-27.5,-176,-24</points>
<connection>
<GID>131</GID>
<name>OUT_2</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-176,-27.5,-172.5,-27.5</points>
<connection>
<GID>184</GID>
<name>IN_2</name></connection>
<intersection>-176 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177,-26.5,-177,-24</points>
<connection>
<GID>131</GID>
<name>OUT_3</name></connection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-177,-26.5,-172.5,-26.5</points>
<connection>
<GID>184</GID>
<name>IN_3</name></connection>
<intersection>-177 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>206.101,21.3898,318.162,-47.6784</PageViewport>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>229,-16.5</position>
<gparam>LABEL_TEXT 4-bit input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>280.5,-16</position>
<gparam>LABEL_TEXT 4-bit input</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>262.5,-26</position>
<gparam>LABEL_TEXT 4-bit output displayed in hex</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>338</ID>
<type>AE_FULLADDER_4BIT</type>
<position>254,-9.5</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>203 </input>
<input>
<ID>IN_2</ID>201 </input>
<input>
<ID>IN_3</ID>199 </input>
<input>
<ID>IN_B_0</ID>185 </input>
<input>
<ID>IN_B_1</ID>186 </input>
<input>
<ID>IN_B_2</ID>187 </input>
<input>
<ID>IN_B_3</ID>188 </input>
<output>
<ID>OUT_0</ID>193 </output>
<output>
<ID>OUT_1</ID>194 </output>
<output>
<ID>OUT_2</ID>195 </output>
<output>
<ID>OUT_3</ID>196 </output>
<input>
<ID>carry_in</ID>197 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>341</ID>
<type>DD_KEYPAD_HEX</type>
<position>225.5,-9</position>
<output>
<ID>OUT_0</ID>204 </output>
<output>
<ID>OUT_1</ID>202 </output>
<output>
<ID>OUT_2</ID>200 </output>
<output>
<ID>OUT_3</ID>198 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>342</ID>
<type>DD_KEYPAD_HEX</type>
<position>276.5,-8</position>
<output>
<ID>OUT_0</ID>185 </output>
<output>
<ID>OUT_1</ID>186 </output>
<output>
<ID>OUT_2</ID>187 </output>
<output>
<ID>OUT_3</ID>188 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>343</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>260,-18</position>
<input>
<ID>IN_0</ID>193 </input>
<input>
<ID>IN_1</ID>194 </input>
<input>
<ID>IN_2</ID>195 </input>
<input>
<ID>IN_3</ID>196 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>345</ID>
<type>EE_VDD</type>
<position>264,-7.5</position>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>347</ID>
<type>AA_LABEL</type>
<position>266,-9.5</position>
<gparam>LABEL_TEXT C_in = 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AE_SMALL_INVERTER</type>
<position>233.5,-5.5</position>
<input>
<ID>IN_0</ID>198 </input>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>351</ID>
<type>AE_SMALL_INVERTER</type>
<position>233.5,-8</position>
<input>
<ID>IN_0</ID>200 </input>
<output>
<ID>OUT_0</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_SMALL_INVERTER</type>
<position>235,-10</position>
<input>
<ID>IN_0</ID>202 </input>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>355</ID>
<type>AE_SMALL_INVERTER</type>
<position>236.5,-12</position>
<input>
<ID>IN_0</ID>204 </input>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_LABEL</type>
<position>226,0.5</position>
<gparam>LABEL_TEXT Input X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>359</ID>
<type>AA_LABEL</type>
<position>279.5,3.5</position>
<gparam>LABEL_TEXT Input Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>361</ID>
<type>AA_LABEL</type>
<position>263,-23</position>
<gparam>LABEL_TEXT Output Z = ?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AA_LABEL</type>
<position>258,12</position>
<gparam>LABEL_TEXT What is the  function Z?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>257.5,8</position>
<gparam>LABEL_TEXT Assume inputs X,Y are 4-bit 2's Complement Nos.</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255.5,-19,255.5,-13.5</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-19,257,-19</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>255.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>254.5,-18,254.5,-13.5</points>
<connection>
<GID>338</GID>
<name>OUT_1</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>254.5,-18,257,-18</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>254.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253.5,-17,253.5,-13.5</points>
<connection>
<GID>338</GID>
<name>OUT_2</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253.5,-17,257,-17</points>
<connection>
<GID>343</GID>
<name>IN_2</name></connection>
<intersection>253.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252.5,-16,252.5,-13.5</points>
<connection>
<GID>338</GID>
<name>OUT_3</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>252.5,-16,257,-16</points>
<connection>
<GID>343</GID>
<name>IN_3</name></connection>
<intersection>252.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>262,-8.5,264,-8.5</points>
<connection>
<GID>345</GID>
<name>OUT_0</name></connection>
<connection>
<GID>338</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-5.5,231.5,-5.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>230.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>230.5,-6,230.5,-5.5</points>
<connection>
<GID>341</GID>
<name>OUT_3</name></connection>
<intersection>-5.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235.5,-5.5,249,-5.5</points>
<connection>
<GID>338</GID>
<name>IN_3</name></connection>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-8,231.5,-8</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<connection>
<GID>341</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-5.5,250,-2.5</points>
<connection>
<GID>338</GID>
<name>IN_2</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>236.5,-2.5,250,-2.5</points>
<intersection>236.5 2</intersection>
<intersection>250 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>236.5,-8,236.5,-2.5</points>
<intersection>-8 3</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>235.5,-8,236.5,-8</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>236.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-10,233,-10</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>341</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>251,-5.5,251,-0.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>238,-0.5,251,-0.5</points>
<intersection>238 2</intersection>
<intersection>251 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>238,-10,238,-0.5</points>
<intersection>-10 3</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>237,-10,238,-10</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>238 2</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>230.5,-12,234.5,-12</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<connection>
<GID>341</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>252,-5.5,252,0.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>239,0.5,252,0.5</points>
<intersection>239 2</intersection>
<intersection>252 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>239,-12,239,0.5</points>
<intersection>-12 3</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>238.5,-12,239,-12</points>
<connection>
<GID>355</GID>
<name>OUT_0</name></connection>
<intersection>239 2</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-5.5,259,0.5</points>
<connection>
<GID>338</GID>
<name>IN_B_0</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,0.5,286,0.5</points>
<intersection>259 0</intersection>
<intersection>286 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>286,-11,286,0.5</points>
<intersection>-11 3</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-11,286,-11</points>
<connection>
<GID>342</GID>
<name>OUT_0</name></connection>
<intersection>286 2</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258,-5.5,258,0</points>
<connection>
<GID>338</GID>
<name>IN_B_1</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>258,0,285,0</points>
<intersection>258 0</intersection>
<intersection>285 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>285,-9,285,0</points>
<intersection>-9 3</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-9,285,-9</points>
<connection>
<GID>342</GID>
<name>OUT_1</name></connection>
<intersection>285 2</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-5.5,257,-0.5</points>
<connection>
<GID>338</GID>
<name>IN_B_2</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-0.5,283.5,-0.5</points>
<intersection>257 0</intersection>
<intersection>283.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>283.5,-7,283.5,-0.5</points>
<intersection>-7 3</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>281.5,-7,283.5,-7</points>
<connection>
<GID>342</GID>
<name>OUT_2</name></connection>
<intersection>283.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>256,-5.5,256,-1</points>
<connection>
<GID>338</GID>
<name>IN_B_3</name></connection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>256,-1,281.5,-1</points>
<intersection>256 0</intersection>
<intersection>281.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>281.5,-5,281.5,-1</points>
<connection>
<GID>342</GID>
<name>OUT_3</name></connection>
<intersection>-1 1</intersection></vsegment></shape></wire></page 4>
<page 5>
<PageViewport>118.02,-72.3622,233.305,-143.418</PageViewport>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>170,-89</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>169.5,-92</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>200,-120</position>
<gparam>LABEL_TEXT =1 if AB=11</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>199.5,-129</position>
<gparam>LABEL_TEXT =0 if AB=00</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>170,-112.5</position>
<gparam>LABEL_TEXT If selectl lines (XY)=10 then Output=Sarah</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>170,-111</position>
<gparam>LABEL_TEXT If selectl lines (XY)=00 then Output= Kevin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>GA_LED</type>
<position>188.5,-120</position>
<input>
<ID>N_in0</ID>179 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>GA_LED</type>
<position>188.5,-123.5</position>
<input>
<ID>N_in0</ID>180 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AE_MUX_4x1</type>
<position>178,-103</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>162 </input>
<input>
<ID>IN_2</ID>163 </input>
<input>
<ID>IN_3</ID>174 </input>
<output>
<ID>OUT</ID>149 </output>
<input>
<ID>SEL_0</ID>154 </input>
<input>
<ID>SEL_1</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>296</ID>
<type>GA_LED</type>
<position>188,-103</position>
<input>
<ID>N_in0</ID>149 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>GA_LED</type>
<position>188.5,-126.5</position>
<input>
<ID>N_in0</ID>181 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>GA_LED</type>
<position>189,-129.5</position>
<input>
<ID>N_in0</ID>182 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>300</ID>
<type>AA_TOGGLE</type>
<position>173,-92</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>301</ID>
<type>EE_VDD</type>
<position>157,-121</position>
<output>
<ID>OUT_0</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>302</ID>
<type>AA_LABEL</type>
<position>172.5,-115</position>
<gparam>LABEL_TEXT Decoder Schematic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>159,-119</position>
<gparam>LABEL_TEXT Voltage source</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>304</ID>
<type>AA_LABEL</type>
<position>162,-123.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>AA_LABEL</type>
<position>162,-126.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>AA_LABEL</type>
<position>168,-129</position>
<gparam>LABEL_TEXT Output selected depends on value of AB</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>AA_LABEL</type>
<position>192.5,-120</position>
<gparam>LABEL_TEXT Linnea</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>308</ID>
<type>AA_LABEL</type>
<position>192,-123</position>
<gparam>LABEL_TEXT Sarah</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>193.5,-126</position>
<gparam>LABEL_TEXT Graham</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>168,-132</position>
<gparam>LABEL_TEXT Output codes go from 0 (00) to 3 (11)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AA_LABEL</type>
<position>192.5,-129</position>
<gparam>LABEL_TEXT Kevin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>AA_LABEL</type>
<position>167,-130.5</position>
<gparam>LABEL_TEXT E is enable signal - enables decoder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_LABEL</type>
<position>170,-133.5</position>
<gparam>LABEL_TEXT Kevin has code 0 (00), Sarah has code 2 (10)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AA_TOGGLE</type>
<position>173,-89</position>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_TOGGLE</type>
<position>164,-99.5</position>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>316</ID>
<type>AA_TOGGLE</type>
<position>164,-102</position>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>317</ID>
<type>AA_TOGGLE</type>
<position>164,-104</position>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_TOGGLE</type>
<position>164,-106</position>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_LABEL</type>
<position>160,-106</position>
<gparam>LABEL_TEXT Kevin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>AA_LABEL</type>
<position>159.5,-104</position>
<gparam>LABEL_TEXT Graham</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>321</ID>
<type>AA_LABEL</type>
<position>160,-102</position>
<gparam>LABEL_TEXT Sarah</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>AA_LABEL</type>
<position>160,-99.5</position>
<gparam>LABEL_TEXT Linnea</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>AA_LABEL</type>
<position>171.5,-85</position>
<gparam>LABEL_TEXT Control Signals (X,Y)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>172.5,-82</position>
<gparam>LABEL_TEXT Multiplexer Schematic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>AA_LABEL</type>
<position>191,-105.5</position>
<gparam>LABEL_TEXT Output</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>AA_LABEL</type>
<position>172.5,-87</position>
<gparam>LABEL_TEXT Determines which input to send to output</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>AA_LABEL</type>
<position>174.5,-109</position>
<gparam>LABEL_TEXT 0 on MUX input lines  indicates this input is select when control signal=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>329</ID>
<type>BA_DECODER_2x4</type>
<position>176.5,-123.5</position>
<input>
<ID>ENABLE</ID>183 </input>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT_0</ID>182 </output>
<output>
<ID>OUT_1</ID>181 </output>
<output>
<ID>OUT_2</ID>180 </output>
<output>
<ID>OUT_3</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AA_TOGGLE</type>
<position>164,-123.5</position>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_TOGGLE</type>
<position>164,-126.5</position>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>181,-103,187,-103</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<connection>
<GID>296</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-98,178,-92</points>
<connection>
<GID>295</GID>
<name>SEL_1</name></connection>
<intersection>-92 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-92,178,-92</points>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection>
<intersection>178 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-98,179,-89</points>
<connection>
<GID>295</GID>
<name>SEL_0</name></connection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-89,179,-89</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-106,175,-106</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-104,175,-104</points>
<connection>
<GID>317</GID>
<name>OUT_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>166,-102,175,-102</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<connection>
<GID>295</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-100,170.5,-99.5</points>
<intersection>-100 2</intersection>
<intersection>-99.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-99.5,170.5,-99.5</points>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170.5,-100,175,-100</points>
<connection>
<GID>295</GID>
<name>IN_3</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-126.5,169.5,-125</points>
<intersection>-126.5 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169.5,-125,173.5,-125</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-126.5,169.5,-126.5</points>
<connection>
<GID>331</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-124,169.5,-123.5</points>
<intersection>-124 2</intersection>
<intersection>-123.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-123.5,169.5,-123.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169.5,-124,173.5,-124</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-122,183.5,-120</points>
<intersection>-122 2</intersection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-120,187.5,-120</points>
<connection>
<GID>293</GID>
<name>N_in0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-122,183.5,-122</points>
<connection>
<GID>329</GID>
<name>OUT_3</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-123.5,183.5,-123</points>
<intersection>-123.5 1</intersection>
<intersection>-123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-123.5,187.5,-123.5</points>
<connection>
<GID>294</GID>
<name>N_in0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-123,183.5,-123</points>
<connection>
<GID>329</GID>
<name>OUT_2</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-126.5,183.5,-124</points>
<intersection>-126.5 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-126.5,187.5,-126.5</points>
<connection>
<GID>297</GID>
<name>N_in0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-124,183.5,-124</points>
<connection>
<GID>329</GID>
<name>OUT_1</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-129.5,183.5,-125</points>
<intersection>-129.5 1</intersection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-129.5,188,-129.5</points>
<connection>
<GID>299</GID>
<name>N_in0</name></connection>
<intersection>183.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179.5,-125,183.5,-125</points>
<connection>
<GID>329</GID>
<name>OUT_0</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>157,-122,173.5,-122</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<connection>
<GID>329</GID>
<name>ENABLE</name></connection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-278.643,224.246,-142.82,140.532</PageViewport>
<gate>
<ID>275</ID>
<type>AA_LABEL</type>
<position>-245,203.5</position>
<gparam>LABEL_TEXT set A=1,B=0,C=1,D=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>276</ID>
<type>AA_MUX_2x1</type>
<position>-233.5,199</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>143 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AA_MUX_2x1</type>
<position>-233.5,192.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>-225.5,196.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_TOGGLE</type>
<position>-240.5,200</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>280</ID>
<type>AA_TOGGLE</type>
<position>-240.5,197.5</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_TOGGLE</type>
<position>-240.5,194</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_TOGGLE</type>
<position>-240.5,190.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_TOGGLE</type>
<position>-238.5,208</position>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>-241,208.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>AA_LABEL</type>
<position>-243,200.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>AA_LABEL</type>
<position>-243,198</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>AA_LABEL</type>
<position>-243,194.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>AA_LABEL</type>
<position>-243,191</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>AA_LABEL</type>
<position>-219,199</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>290</ID>
<type>GA_LED</type>
<position>-218,196.5</position>
<input>
<ID>N_in0</ID>148 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>291</ID>
<type>AA_LABEL</type>
<position>-233.5,213</position>
<gparam>LABEL_TEXT What is the function F ?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_LABEL</type>
<position>-230.5,210.5</position>
<gparam>LABEL_TEXT (for x=0? for x=1?)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>-233.5,187.5</position>
<gparam>LABEL_TEXT MUX notation: Input at line 0 is selected if x=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,197.5,-230,199</points>
<intersection>197.5 1</intersection>
<intersection>199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230,197.5,-228.5,197.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>-230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-231.5,199,-230,199</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>-230 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,192.5,-230,195.5</points>
<intersection>192.5 2</intersection>
<intersection>195.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230,195.5,-228.5,195.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>-230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-231.5,192.5,-230,192.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>-230 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-238.5,200,-235.5,200</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<connection>
<GID>276</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237,197.5,-237,198</points>
<intersection>197.5 2</intersection>
<intersection>198 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-237,198,-235.5,198</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>-237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-238.5,197.5,-237,197.5</points>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>-237 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237,193.5,-237,194</points>
<intersection>193.5 1</intersection>
<intersection>194 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-237,193.5,-235.5,193.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>-237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-238.5,194,-237,194</points>
<connection>
<GID>281</GID>
<name>OUT_0</name></connection>
<intersection>-237 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237,190.5,-237,191.5</points>
<intersection>190.5 2</intersection>
<intersection>191.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-237,191.5,-235.5,191.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>-237 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-238.5,190.5,-237,190.5</points>
<connection>
<GID>282</GID>
<name>OUT_0</name></connection>
<intersection>-237 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-231,195,-231,208</points>
<intersection>195 2</intersection>
<intersection>201.5 3</intersection>
<intersection>208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-236.5,208,-231,208</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>-231 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,195,-231,195</points>
<connection>
<GID>277</GID>
<name>SEL_0</name></connection>
<intersection>-231 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-233.5,201.5,-231,201.5</points>
<connection>
<GID>276</GID>
<name>SEL_0</name></connection>
<intersection>-231 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-222.5,196.5,-219,196.5</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>290</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>71.5912,-134.242,194.934,-210.264</PageViewport>
<gate>
<ID>193</ID>
<type>AA_MUX_2x1</type>
<position>132.5,-198.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>209 </input>
<output>
<ID>OUT</ID>192 </output>
<input>
<ID>SEL_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>169.5,-180</position>
<gparam>LABEL_TEXT 4-bit Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>122.5,-154.5</position>
<output>
<ID>OUT_0</ID>136 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>123.5,-151.5</position>
<gparam>LABEL_TEXT Input C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>170.5,-191</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>140 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 13</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_FULLADDER_4BIT</type>
<position>157,-179.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>206 </input>
<input>
<ID>IN_2</ID>207 </input>
<input>
<ID>IN_3</ID>208 </input>
<input>
<ID>IN_B_0</ID>184 </input>
<input>
<ID>IN_B_1</ID>189 </input>
<input>
<ID>IN_B_2</ID>190 </input>
<input>
<ID>IN_B_3</ID>191 </input>
<output>
<ID>OUT_0</ID>137 </output>
<output>
<ID>OUT_1</ID>138 </output>
<output>
<ID>OUT_2</ID>139 </output>
<output>
<ID>OUT_3</ID>140 </output>
<input>
<ID>carry_in</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>205</ID>
<type>AE_SMALL_INVERTER</type>
<position>127.5,-197.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>123,-191.5</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>120,-185.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>137</ID>
<type>AE_SMALL_INVERTER</type>
<position>118,-179.5</position>
<input>
<ID>IN_0</ID>135 </input>
<output>
<ID>OUT_0</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>133,-144.5</position>
<gparam>LABEL_TEXT Describe what this circuit/device does? </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>128,-147.5</position>
<gparam>LABEL_TEXT Inputs: X,Y,C and Output: F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>DD_KEYPAD_HEX</type>
<position>103,-164</position>
<output>
<ID>OUT_0</ID>184 </output>
<output>
<ID>OUT_1</ID>189 </output>
<output>
<ID>OUT_2</ID>190 </output>
<output>
<ID>OUT_3</ID>191 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>168.5,-196</position>
<gparam>LABEL_TEXT 4-bit output F</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>148.5,-150.5</position>
<gparam>LABEL_TEXT X,Y are 4-bit 2s complement numbers</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>DD_KEYPAD_HEX</type>
<position>103.5,-194.5</position>
<output>
<ID>OUT_0</ID>123 </output>
<output>
<ID>OUT_1</ID>124 </output>
<output>
<ID>OUT_2</ID>134 </output>
<output>
<ID>OUT_3</ID>135 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 6</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>96,-170</position>
<gparam>LABEL_TEXT Input Y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_LABEL</type>
<position>95.5,-193</position>
<gparam>LABEL_TEXT Input X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_MUX_2x1</type>
<position>128,-192.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>206 </output>
<input>
<ID>SEL_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_MUX_2x1</type>
<position>125,-186.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>207 </output>
<input>
<ID>SEL_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_MUX_2x1</type>
<position>122.5,-180.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>208 </output>
<input>
<ID>SEL_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-175.5,154,-172</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-172 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-172,154,-172</points>
<intersection>130 2</intersection>
<intersection>154 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>130,-192.5,130,-172</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>-172 1</intersection></vsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153,-175.5,153,-173</points>
<connection>
<GID>203</GID>
<name>IN_2</name></connection>
<intersection>-173 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-173,153,-173</points>
<intersection>127 2</intersection>
<intersection>153 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>127,-186.5,127,-173</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>-173 1</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-175.5,152,-174</points>
<connection>
<GID>203</GID>
<name>IN_3</name></connection>
<intersection>-174 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-174,152,-174</points>
<intersection>124.5 2</intersection>
<intersection>152 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>124.5,-180.5,124.5,-174</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>-174 1</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129.5,-197.5,130.5,-197.5</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<connection>
<GID>193</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-191.5,126,-191.5</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<connection>
<GID>185</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122,-185.5,123,-185.5</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,-179.5,120.5,-179.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<connection>
<GID>189</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>108.5,-197.5,125.5,-197.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>108.5 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>108.5,-199.5,108.5,-197.5</points>
<intersection>-199.5 16</intersection>
<intersection>-197.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>108.5,-199.5,130.5,-199.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>108.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-195.5,117.5,-193.5</points>
<intersection>-195.5 2</intersection>
<intersection>-193.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117.5,-193.5,126,-193.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>117.5 0</intersection>
<intersection>121 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-195.5,117.5,-195.5</points>
<connection>
<GID>151</GID>
<name>OUT_1</name></connection>
<intersection>117.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121,-193.5,121,-191.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>-193.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-193.5,115.5,-187.5</points>
<intersection>-193.5 2</intersection>
<intersection>-187.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-187.5,123,-187.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection>
<intersection>118 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-193.5,115.5,-193.5</points>
<connection>
<GID>151</GID>
<name>OUT_2</name></connection>
<intersection>115.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118,-187.5,118,-185.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-187.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-191.5,114.5,-181.5</points>
<intersection>-191.5 2</intersection>
<intersection>-181.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-181.5,120.5,-181.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection>
<intersection>116 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>108.5,-191.5,114.5,-191.5</points>
<connection>
<GID>151</GID>
<name>OUT_3</name></connection>
<intersection>114.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>116,-181.5,116,-179.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-181.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124.5,-154.5,165,-154.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>132.5 2</intersection>
<intersection>165 10</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>132.5,-196,132.5,-154.5</points>
<connection>
<GID>193</GID>
<name>SEL_0</name></connection>
<intersection>-188 5</intersection>
<intersection>-184 6</intersection>
<intersection>-178 4</intersection>
<intersection>-154.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>122.5,-178,132.5,-178</points>
<connection>
<GID>189</GID>
<name>SEL_0</name></connection>
<intersection>132.5 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>128,-188,132.5,-188</points>
<intersection>128 8</intersection>
<intersection>132.5 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>125,-184,132.5,-184</points>
<connection>
<GID>187</GID>
<name>SEL_0</name></connection>
<intersection>132.5 2</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>128,-190,128,-188</points>
<connection>
<GID>185</GID>
<name>SEL_0</name></connection>
<intersection>-188 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>165,-178.5,165,-154.5</points>
<connection>
<GID>203</GID>
<name>carry_in</name></connection>
<intersection>-154.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>158.5,-192,158.5,-183.5</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<intersection>-192 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158.5,-192,167.5,-192</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>158.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157.5,-191,157.5,-183.5</points>
<connection>
<GID>203</GID>
<name>OUT_1</name></connection>
<intersection>-191 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157.5,-191,167.5,-191</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>157.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-190,156.5,-183.5</points>
<connection>
<GID>203</GID>
<name>OUT_2</name></connection>
<intersection>-190 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-190,167.5,-190</points>
<connection>
<GID>201</GID>
<name>IN_2</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-189,155.5,-183.5</points>
<connection>
<GID>203</GID>
<name>OUT_3</name></connection>
<intersection>-189 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155.5,-189,167.5,-189</points>
<connection>
<GID>201</GID>
<name>IN_3</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-175.5,162,-167</points>
<connection>
<GID>203</GID>
<name>IN_B_0</name></connection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-167,162,-167</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>162 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-175.5,161,-165</points>
<connection>
<GID>203</GID>
<name>IN_B_1</name></connection>
<intersection>-165 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-165,161,-165</points>
<connection>
<GID>142</GID>
<name>OUT_1</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-175.5,160,-163</points>
<connection>
<GID>203</GID>
<name>IN_B_2</name></connection>
<intersection>-163 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-163,160,-163</points>
<connection>
<GID>142</GID>
<name>OUT_2</name></connection>
<intersection>160 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-175.5,159,-161</points>
<connection>
<GID>203</GID>
<name>IN_B_3</name></connection>
<intersection>-161 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-161,159,-161</points>
<connection>
<GID>142</GID>
<name>OUT_3</name></connection>
<intersection>159 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143.5,-198.5,143.5,-171</points>
<intersection>-198.5 1</intersection>
<intersection>-171 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134.5,-198.5,143.5,-198.5</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<intersection>143.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143.5,-171,155,-171</points>
<intersection>143.5 0</intersection>
<intersection>155 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>155,-175.5,155,-171</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-171 2</intersection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>-96.8735,171.766,-7.97649,116.975</PageViewport>
<gate>
<ID>207</ID>
<type>AA_MUX_2x1</type>
<position>-67,145.5</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>254 </input>
<output>
<ID>OUT</ID>240 </output>
<input>
<ID>SEL_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_MUX_2x1</type>
<position>-63.5,138.5</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>241 </output>
<input>
<ID>SEL_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_MUX_2x1</type>
<position>-59,131</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>242 </output>
<input>
<ID>SEL_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_MUX_2x1</type>
<position>-55,123.5</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>243 </output>
<input>
<ID>SEL_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>BA_DECODER_2x4</type>
<position>-76,164</position>
<input>
<ID>ENABLE</ID>229 </input>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT_0</ID>245 </output>
<output>
<ID>OUT_1</ID>246 </output>
<output>
<ID>OUT_2</ID>247 </output>
<output>
<ID>OUT_3</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>-71,144.5</position>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>-68,137.5</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>-63.5,128.5</position>
<output>
<ID>OUT_0</ID>251 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>-60.5,122.5</position>
<output>
<ID>OUT_0</ID>252 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>-72.5,144.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>-70,137.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>-65.5,129.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>-62,122</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_TOGGLE</type>
<position>-81,153.5</position>
<output>
<ID>OUT_0</ID>253 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>-81,150</position>
<output>
<ID>OUT_0</ID>244 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_AND2</type>
<position>-74.5,151.5</position>
<input>
<ID>IN_0</ID>253 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_TOGGLE</type>
<position>-81,139.5</position>
<output>
<ID>OUT_0</ID>232 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_TOGGLE</type>
<position>-81,129.5</position>
<output>
<ID>OUT_0</ID>235 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>-80.5,124.5</position>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_TOGGLE</type>
<position>-80.5,119.5</position>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_TOGGLE</type>
<position>-86,163</position>
<output>
<ID>OUT_0</ID>256 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_TOGGLE</type>
<position>-86,160</position>
<output>
<ID>OUT_0</ID>255 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>-88,163</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>273</ID>
<type>AA_LABEL</type>
<position>-88,160</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>AA_LABEL</type>
<position>-84,153.5</position>
<gparam>LABEL_TEXT x0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>AA_LABEL</type>
<position>-84,150</position>
<gparam>LABEL_TEXT y0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>333</ID>
<type>AA_LABEL</type>
<position>-85.5,143</position>
<gparam>LABEL_TEXT x1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>334</ID>
<type>AA_LABEL</type>
<position>-85,130.5</position>
<gparam>LABEL_TEXT y2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>335</ID>
<type>AA_LABEL</type>
<position>-84,124.5</position>
<gparam>LABEL_TEXT x3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>336</ID>
<type>AA_LABEL</type>
<position>-84,119.5</position>
<gparam>LABEL_TEXT y3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>GA_LED</type>
<position>-33,142</position>
<input>
<ID>N_in0</ID>239 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>339</ID>
<type>AA_AND2</type>
<position>-71.5,123.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_TOGGLE</type>
<position>-81.5,142.5</position>
<output>
<ID>OUT_0</ID>231 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_TOGGLE</type>
<position>-81,133</position>
<output>
<ID>OUT_0</ID>234 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>346</ID>
<type>AA_LABEL</type>
<position>-85,139.5</position>
<gparam>LABEL_TEXT y1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>348</ID>
<type>AA_LABEL</type>
<position>-84.5,133.5</position>
<gparam>LABEL_TEXT x2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>350</ID>
<type>AE_OR4</type>
<position>-42,142.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<input>
<ID>IN_2</ID>242 </input>
<input>
<ID>IN_3</ID>243 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_LABEL</type>
<position>-75.5,160.5</position>
<gparam>LABEL_TEXT 4-1 decoder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>-54,118</position>
<gparam>LABEL_TEXT 2-1 MUX</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>356</ID>
<type>AA_LABEL</type>
<position>-49,171</position>
<gparam>LABEL_TEXT What is the function F computed by circuit?</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>AA_LABEL</type>
<position>-33,146</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>360</ID>
<type>AA_LABEL</type>
<position>-33.5,155.5</position>
<gparam>LABEL_TEXT which output from decoder is enabled?</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>AA_LABEL</type>
<position>-33,153.5</position>
<gparam>LABEL_TEXT which multiplexer will have select line=1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>364</ID>
<type>AA_AND2</type>
<position>-73.5,140.5</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AA_AND2</type>
<position>-69.5,132</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>-41,164.5</position>
<gparam>LABEL_TEXT Input to decoder: A,B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>368</ID>
<type>EE_VDD</type>
<position>-82.5,166.5</position>
<output>
<ID>OUT_0</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_LABEL</type>
<position>-38,162</position>
<gparam>LABEL_TEXT Other inputs: x0,..,x3,y0..,y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>AA_LABEL</type>
<position>-45.5,160</position>
<gparam>LABEL_TEXT Output= F</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>371</ID>
<type>AA_LABEL</type>
<position>-36.5,157.5</position>
<gparam>LABEL_TEXT Hint: If A=0,B=0 what is output function F</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82.5,165.5,-79,165.5</points>
<connection>
<GID>368</GID>
<name>OUT_0</name></connection>
<connection>
<GID>243</GID>
<name>ENABLE</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,139.5,-68,140.5</points>
<intersection>139.5 1</intersection>
<intersection>140.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,139.5,-65.5,139.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>-68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,140.5,-68,140.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,141.5,-78,142.5</points>
<intersection>141.5 1</intersection>
<intersection>142.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,141.5,-76.5,141.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,142.5,-78,142.5</points>
<connection>
<GID>340</GID>
<name>OUT_0</name></connection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,139.5,-76.5,139.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<connection>
<GID>364</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66.5,132,-61,132</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<connection>
<GID>366</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,133,-72.5,133</points>
<connection>
<GID>344</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76,129.5,-76,131</points>
<intersection>129.5 2</intersection>
<intersection>131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,131,-72.5,131</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>-76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,129.5,-76,129.5</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>-76 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,123.5,-63,124.5</points>
<intersection>123.5 2</intersection>
<intersection>124.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,124.5,-57,124.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,123.5,-63,123.5</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-78.5,124.5,-74.5,124.5</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,119.5,-76.5,122.5</points>
<intersection>119.5 2</intersection>
<intersection>122.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,122.5,-74.5,122.5</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,119.5,-76.5,119.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38,142.5,-34,142.5</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<intersection>-34 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-34,142,-34,142.5</points>
<connection>
<GID>337</GID>
<name>N_in0</name></connection>
<intersection>142.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-65,145.5,-45,145.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<connection>
<GID>350</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,138.5,-53.5,143.5</points>
<intersection>138.5 2</intersection>
<intersection>143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53.5,143.5,-45,143.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-61.5,138.5,-53.5,138.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,131,-51,141.5</points>
<intersection>131 1</intersection>
<intersection>141.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57,131,-51,131</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>-51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-51,141.5,-45,141.5</points>
<connection>
<GID>350</GID>
<name>IN_2</name></connection>
<intersection>-51 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,123.5,-49,139.5</points>
<intersection>123.5 1</intersection>
<intersection>139.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-53,123.5,-49,123.5</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>-49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-49,139.5,-45,139.5</points>
<connection>
<GID>350</GID>
<name>IN_3</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,150,-78.5,150.5</points>
<intersection>150 1</intersection>
<intersection>150.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-79,150,-78.5,150</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-78.5,150.5,-77.5,150.5</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67,148,-67,162.5</points>
<connection>
<GID>207</GID>
<name>SEL_0</name></connection>
<intersection>162.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,162.5,-67,162.5</points>
<connection>
<GID>243</GID>
<name>OUT_0</name></connection>
<intersection>-67 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,141,-63.5,163.5</points>
<connection>
<GID>225</GID>
<name>SEL_0</name></connection>
<intersection>163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,163.5,-63.5,163.5</points>
<connection>
<GID>243</GID>
<name>OUT_1</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59,133.5,-59,164.5</points>
<connection>
<GID>231</GID>
<name>SEL_0</name></connection>
<intersection>164.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,164.5,-59,164.5</points>
<connection>
<GID>243</GID>
<name>OUT_2</name></connection>
<intersection>-59 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,126,-55,165.5</points>
<connection>
<GID>232</GID>
<name>SEL_0</name></connection>
<intersection>165.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,165.5,-55,165.5</points>
<connection>
<GID>243</GID>
<name>OUT_3</name></connection>
<intersection>-55 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-69,144.5,-69,144.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66,137.5,-65.5,137.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-61,128.5,-61,130</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>128.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-61.5,128.5,-61,128.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-61 2</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58.5,122.5,-57,122.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,152.5,-78.5,153.5</points>
<intersection>152.5 1</intersection>
<intersection>153.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78.5,152.5,-77.5,152.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,153.5,-78.5,153.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>-78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,146.5,-70.5,151.5</points>
<intersection>146.5 1</intersection>
<intersection>151.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-70.5,146.5,-69,146.5</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>-70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,151.5,-70.5,151.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,160,-81.5,162.5</points>
<intersection>160 2</intersection>
<intersection>162.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81.5,162.5,-79,162.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-84,160,-81.5,160</points>
<connection>
<GID>271</GID>
<name>OUT_0</name></connection>
<intersection>-81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,163,-81.5,163.5</points>
<intersection>163 2</intersection>
<intersection>163.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-81.5,163.5,-79,163.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-84,163,-81.5,163</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>-81.5 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>304.099,15.0909,544.505,-133.083</PageViewport>
<gate>
<ID>266</ID>
<type>FF_GND</type>
<position>429,-30.5</position>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>447.5,-16.5</position>
<gparam>LABEL_TEXT Input C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>456.5,-20</position>
<gparam>LABEL_TEXT (control signal)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>391.5,-75.5</position>
<gparam>LABEL_TEXT Comparator: one of three outputs is a 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>391.5,-84</position>
<gparam>LABEL_TEXT (output=1 if X>Y, 2 if X=Y, 4 if XY )</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AE_FULLADDER_4BIT</type>
<position>414.5,-23</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>88 </input>
<input>
<ID>IN_2</ID>87 </input>
<input>
<ID>IN_3</ID>86 </input>
<input>
<ID>IN_B_0</ID>85 </input>
<input>
<ID>IN_B_1</ID>84 </input>
<input>
<ID>IN_B_2</ID>82 </input>
<input>
<ID>IN_B_3</ID>81 </input>
<output>
<ID>OUT_0</ID>105 </output>
<output>
<ID>OUT_1</ID>106 </output>
<output>
<ID>OUT_2</ID>107 </output>
<output>
<ID>OUT_3</ID>108 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>158</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>416,-60</position>
<output>
<ID>A_equal_B</ID>103 </output>
<output>
<ID>A_greater_B</ID>102 </output>
<output>
<ID>A_less_B</ID>104 </output>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>97 </input>
<input>
<ID>IN_B_0</ID>93 </input>
<input>
<ID>IN_B_1</ID>92 </input>
<input>
<ID>IN_B_2</ID>91 </input>
<input>
<ID>IN_B_3</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>337.5,-2.5</position>
<gparam>LABEL_TEXT Number Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>339,-74.5</position>
<gparam>LABEL_TEXT Number X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>412.5,-12</position>
<gparam>LABEL_TEXT Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_MUX_2x1</type>
<position>433,-26.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>101 </output>
<input>
<ID>SEL_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_MUX_2x1</type>
<position>433,-35.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>100 </output>
<input>
<ID>SEL_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_MUX_2x1</type>
<position>433,-44.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>99 </output>
<input>
<ID>SEL_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_MUX_2x1</type>
<position>433,-54</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>98 </output>
<input>
<ID>SEL_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>455.5,-41</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>99 </input>
<input>
<ID>IN_2</ID>100 </input>
<input>
<ID>IN_3</ID>101 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>442,-20.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>373.5,7.5</position>
<gparam>LABEL_TEXT What does this circuit do..</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>HE_JUNC_4</type>
<position>373.5,-9</position>
<input>
<ID>N_in0</ID>74 </input>
<input>
<ID>N_in1</ID>81 </input>
<input>
<ID>N_in2</ID>90 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>HE_JUNC_4</type>
<position>375,-11</position>
<input>
<ID>N_in0</ID>75 </input>
<input>
<ID>N_in1</ID>82 </input>
<input>
<ID>N_in2</ID>91 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>HE_JUNC_4</type>
<position>378,-15</position>
<input>
<ID>N_in0</ID>76 </input>
<input>
<ID>N_in1</ID>85 </input>
<input>
<ID>N_in2</ID>93 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>HE_JUNC_4</type>
<position>359,-56</position>
<input>
<ID>N_in0</ID>77 </input>
<input>
<ID>N_in2</ID>97 </input>
<input>
<ID>N_in3</ID>86 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>HE_JUNC_4</type>
<position>361.5,-58</position>
<input>
<ID>N_in0</ID>78 </input>
<input>
<ID>N_in2</ID>96 </input>
<input>
<ID>N_in3</ID>87 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>HE_JUNC_4</type>
<position>365,-60</position>
<input>
<ID>N_in0</ID>79 </input>
<input>
<ID>N_in2</ID>95 </input>
<input>
<ID>N_in3</ID>88 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>HE_JUNC_4</type>
<position>368,-62</position>
<input>
<ID>N_in0</ID>80 </input>
<input>
<ID>N_in1</ID>94 </input>
<input>
<ID>N_in3</ID>89 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>DD_KEYPAD_HEX</type>
<position>350,-59</position>
<output>
<ID>OUT_0</ID>80 </output>
<output>
<ID>OUT_1</ID>79 </output>
<output>
<ID>OUT_2</ID>78 </output>
<output>
<ID>OUT_3</ID>77 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>177</ID>
<type>HE_JUNC_4</type>
<position>376.5,-13</position>
<input>
<ID>N_in0</ID>83 </input>
<input>
<ID>N_in1</ID>84 </input>
<input>
<ID>N_in2</ID>92 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>DD_KEYPAD_HEX</type>
<position>349.5,-12</position>
<output>
<ID>OUT_0</ID>76 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>75 </output>
<output>
<ID>OUT_3</ID>74 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>392,-81.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>436.5,-57.5</position>
<gparam>LABEL_TEXT 2-1 Multiplexer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>AA_LABEL</type>
<position>392,-80</position>
<gparam>LABEL_TEXT Signal at > is 1 if X>Y, E is 1 if equal,  is 1 if XY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-9,372.5,-9</points>
<connection>
<GID>178</GID>
<name>OUT_3</name></connection>
<connection>
<GID>169</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-11,374,-11</points>
<connection>
<GID>178</GID>
<name>OUT_2</name></connection>
<connection>
<GID>170</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-15,377,-15</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<connection>
<GID>171</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,-56,358,-56</points>
<connection>
<GID>176</GID>
<name>OUT_3</name></connection>
<connection>
<GID>172</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,-58,360.5,-58</points>
<connection>
<GID>176</GID>
<name>OUT_2</name></connection>
<connection>
<GID>173</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,-60,364,-60</points>
<connection>
<GID>176</GID>
<name>OUT_1</name></connection>
<connection>
<GID>174</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>355,-62,367,-62</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<connection>
<GID>175</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>385,-21,385,-9</points>
<intersection>-21 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>385,-21,410.5,-21</points>
<connection>
<GID>157</GID>
<name>IN_B_3</name></connection>
<intersection>385 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>374.5,-9,385,-9</points>
<connection>
<GID>169</GID>
<name>N_in1</name></connection>
<intersection>385 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386,-20,386,-11</points>
<intersection>-20 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>386,-20,410.5,-20</points>
<connection>
<GID>157</GID>
<name>IN_B_2</name></connection>
<intersection>386 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>376,-11,386,-11</points>
<connection>
<GID>170</GID>
<name>N_in1</name></connection>
<intersection>386 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-13,375.5,-13</points>
<connection>
<GID>178</GID>
<name>OUT_1</name></connection>
<connection>
<GID>177</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>388,-19,388,-13</points>
<intersection>-19 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>388,-19,410.5,-19</points>
<connection>
<GID>157</GID>
<name>IN_B_1</name></connection>
<intersection>388 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>377.5,-13,388,-13</points>
<connection>
<GID>177</GID>
<name>N_in1</name></connection>
<intersection>388 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389.5,-18,389.5,-15</points>
<intersection>-18 1</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>389.5,-18,410.5,-18</points>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection>
<intersection>389.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>379,-15,389.5,-15</points>
<connection>
<GID>171</GID>
<name>N_in1</name></connection>
<intersection>389.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-55,359,-28</points>
<connection>
<GID>172</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-28,410.5,-28</points>
<connection>
<GID>157</GID>
<name>IN_3</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-57,361.5,-27</points>
<connection>
<GID>173</GID>
<name>N_in3</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-27,410.5,-27</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365,-59,365,-26</points>
<connection>
<GID>174</GID>
<name>N_in3</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365,-26,410.5,-26</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>365 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>368,-61,368,-25</points>
<connection>
<GID>175</GID>
<name>N_in3</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>368,-25,410.5,-25</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>368 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373.5,-58,373.5,-10</points>
<connection>
<GID>169</GID>
<name>N_in2</name></connection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373.5,-58,412,-58</points>
<connection>
<GID>158</GID>
<name>IN_B_3</name></connection>
<intersection>373.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>375,-57,375,-12</points>
<connection>
<GID>170</GID>
<name>N_in2</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>375,-57,412,-57</points>
<connection>
<GID>158</GID>
<name>IN_B_2</name></connection>
<intersection>375 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376.5,-56,376.5,-14</points>
<connection>
<GID>177</GID>
<name>N_in2</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>376.5,-56,412,-56</points>
<connection>
<GID>158</GID>
<name>IN_B_1</name></connection>
<intersection>376.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>378,-55,378,-16</points>
<connection>
<GID>171</GID>
<name>N_in2</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>378,-55,412,-55</points>
<connection>
<GID>158</GID>
<name>IN_B_0</name></connection>
<intersection>378 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>369,-62,412,-62</points>
<connection>
<GID>175</GID>
<name>N_in1</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>365,-63.5,365,-61</points>
<connection>
<GID>174</GID>
<name>N_in2</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365,-63.5,412,-63.5</points>
<intersection>365 0</intersection>
<intersection>412 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>412,-63.5,412,-63</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>-63.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>361.5,-64,361.5,-59</points>
<connection>
<GID>173</GID>
<name>N_in2</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>361.5,-64,412,-64</points>
<connection>
<GID>158</GID>
<name>IN_2</name></connection>
<intersection>361.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-65,359,-57</points>
<connection>
<GID>172</GID>
<name>N_in2</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-65,412,-65</points>
<connection>
<GID>158</GID>
<name>IN_3</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>444.5,-54,444.5,-42</points>
<intersection>-54 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435,-54,444.5,-54</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>444.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>444.5,-42,452.5,-42</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>444.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443.5,-44.5,443.5,-41</points>
<intersection>-44.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435,-44.5,443.5,-44.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443.5,-41,452.5,-41</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>443.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>443.5,-40,443.5,-35.5</points>
<intersection>-40 2</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435,-35.5,443.5,-35.5</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>443.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>443.5,-40,452.5,-40</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>443.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>446,-39,446,-26.5</points>
<intersection>-39 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>435,-26.5,446,-26.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>446 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>446,-39,452.5,-39</points>
<connection>
<GID>166</GID>
<name>IN_3</name></connection>
<intersection>446 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>414,-73.5,414,-68</points>
<connection>
<GID>158</GID>
<name>A_greater_B</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>414,-73.5,431,-73.5</points>
<intersection>414 0</intersection>
<intersection>431 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>431,-73.5,431,-55</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>416,-72.5,416,-68</points>
<connection>
<GID>158</GID>
<name>A_equal_B</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>416,-72.5,428.5,-72.5</points>
<intersection>416 0</intersection>
<intersection>428.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>428.5,-72.5,428.5,-45.5</points>
<intersection>-72.5 1</intersection>
<intersection>-45.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>428.5,-45.5,431,-45.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>428.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>426.5,-68,426.5,-36.5</points>
<intersection>-68 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>426.5,-36.5,431,-36.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>426.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>418,-68,426.5,-68</points>
<connection>
<GID>158</GID>
<name>A_less_B</name></connection>
<intersection>426.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421,-53,421,-21.5</points>
<intersection>-53 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418.5,-21.5,421,-21.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>421 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421,-53,431,-53</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>421 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>422.5,-43.5,422.5,-22.5</points>
<intersection>-43.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418.5,-22.5,422.5,-22.5</points>
<connection>
<GID>157</GID>
<name>OUT_1</name></connection>
<intersection>422.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>422.5,-43.5,431,-43.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>422.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-34.5,423.5,-23.5</points>
<intersection>-34.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418.5,-23.5,423.5,-23.5</points>
<connection>
<GID>157</GID>
<name>OUT_2</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>423.5,-34.5,431,-34.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-25.5,424.5,-24.5</points>
<intersection>-25.5 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>418.5,-24.5,424.5,-24.5</points>
<connection>
<GID>157</GID>
<name>OUT_3</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>424.5,-25.5,431,-25.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>437,-51.5,437,-20.5</points>
<intersection>-51.5 8</intersection>
<intersection>-42 9</intersection>
<intersection>-33 10</intersection>
<intersection>-24 11</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>437,-20.5,440,-20.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>433,-51.5,437,-51.5</points>
<connection>
<GID>165</GID>
<name>SEL_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>433,-42,437,-42</points>
<connection>
<GID>164</GID>
<name>SEL_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>433,-33,437,-33</points>
<connection>
<GID>163</GID>
<name>SEL_0</name></connection>
<intersection>437 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>433,-24,437,-24</points>
<connection>
<GID>162</GID>
<name>SEL_0</name></connection>
<intersection>437 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429,-29.5,429,-27.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429,-27.5,431,-27.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>429 0</intersection></hsegment></shape></wire></page 9></circuit>