<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>315.578,-182.734,403.512,-234.014</PageViewport>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW_NT</type>
<position>356,-242.5</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUTINV_0</ID>4 </output>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>355,-231</position>
<gparam>LABEL_TEXT D Flip Flop Schematic</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>331,-240.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>BB_CLOCK</type>
<position>332.5,-252.5</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>371.5,-240.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>350,-199.5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>363,-193</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>365,-205.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>BA_NAND2</type>
<position>368,-195.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>368.5,-203.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>HA_JUNC_2</type>
<position>360.5,-194.5</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>5 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>HA_JUNC_2</type>
<position>360.5,-204.5</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>6 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>HE_JUNC_4</type>
<position>373,-203.5</position>
<input>
<ID>N_in0</ID>7 </input>
<input>
<ID>N_in3</ID>8 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>HE_JUNC_4</type>
<position>373.5,-195.5</position>
<input>
<ID>N_in0</ID>9 </input>
<input>
<ID>N_in1</ID>40 </input>
<input>
<ID>N_in2</ID>10 </input>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>333,-193.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>338.5,-190.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>BA_NAND2</type>
<position>350.5,-195</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND2</type>
<position>350.5,-205</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>341,-206</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>HE_JUNC_4</type>
<position>339,-193.5</position>
<input>
<ID>N_in0</ID>13 </input>
<input>
<ID>N_in1</ID>12 </input>
<input>
<ID>N_in2</ID>14 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>HE_JUNC_4</type>
<position>347,-200</position>
<input>
<ID>N_in2</ID>38 </input>
<input>
<ID>N_in3</ID>15 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>395.5,-201</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>409,-194.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>411,-207</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>BA_NAND2</type>
<position>414,-197</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>414.5,-205</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>HA_JUNC_2</type>
<position>406.5,-196</position>
<input>
<ID>N_in0</ID>36 </input>
<input>
<ID>N_in1</ID>18 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>HA_JUNC_2</type>
<position>406.5,-206</position>
<input>
<ID>N_in0</ID>37 </input>
<input>
<ID>N_in1</ID>19 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>HE_JUNC_4</type>
<position>419,-205</position>
<input>
<ID>N_in0</ID>20 </input>
<input>
<ID>N_in3</ID>21 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>HE_JUNC_4</type>
<position>419.5,-197</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>24 </input>
<input>
<ID>N_in2</ID>23 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>425.5,-197</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>392,-193</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>BA_NAND2</type>
<position>396.5,-196.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>BA_NAND2</type>
<position>396.5,-206.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AE_SMALL_INVERTER</type>
<position>391,-207.5</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>42</ID>
<type>HE_JUNC_4</type>
<position>391,-195.5</position>
<input>
<ID>N_in0</ID>40 </input>
<input>
<ID>N_in1</ID>32 </input>
<input>
<ID>N_in2</ID>33 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>HE_JUNC_4</type>
<position>393,-201.5</position>
<input>
<ID>N_in0</ID>39 </input>
<input>
<ID>N_in2</ID>35 </input>
<input>
<ID>N_in3</ID>34 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AE_SMALL_INVERTER</type>
<position>363.5,-216</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>BB_CLOCK</type>
<position>366.5,-220.5</position>
<output>
<ID>CLK</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>373.5,-190.5</position>
<input>
<ID>N_in2</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>380,-188</position>
<gparam>LABEL_TEXT Q_intermediate</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>427,-192.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>370,-183.5</position>
<gparam>LABEL_TEXT D Flip-Flop</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>325.5,-237</position>
<gparam>LABEL_TEXT Input D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>326,-248</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>366.5,-237.5</position>
<gparam>LABEL_TEXT Output Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>368.5,-248</position>
<gparam>LABEL_TEXT Output Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>371,-244</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>406.5,-231</position>
<gparam>LABEL_TEXT D Flip-flop with write enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AF_DFF_LOW</type>
<position>406,-244</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>50 </input>
<input>
<ID>clock_enable</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>397,-240.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_TOGGLE</type>
<position>396,-247</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>413.5,-241.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>BB_CLOCK</type>
<position>389.5,-243.5</position>
<output>
<ID>CLK</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>344.5,-252.5,344.5,-243.5</points>
<intersection>-252.5 2</intersection>
<intersection>-243.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>344.5,-243.5,353,-243.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>344.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>336.5,-252.5,344.5,-252.5</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<intersection>344.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>333,-240.5,353,-240.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>359,-240.5,370.5,-240.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>370.5,-244,370.5,-243.5</points>
<intersection>-244 1</intersection>
<intersection>-243.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>370,-244,370.5,-244</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<intersection>370.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>359,-243.5,370.5,-243.5</points>
<connection>
<GID>1</GID>
<name>OUTINV_0</name></connection>
<intersection>370.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361.5,-194.5,365,-194.5</points>
<connection>
<GID>11</GID>
<name>N_in1</name></connection>
<connection>
<GID>9</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>361.5,-204.5,365.5,-204.5</points>
<connection>
<GID>12</GID>
<name>N_in1</name></connection>
<connection>
<GID>10</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>371.5,-203.5,372,-203.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<connection>
<GID>13</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,-202.5,373,-199</points>
<connection>
<GID>13</GID>
<name>N_in3</name></connection>
<intersection>-199 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>365,-199,373,-199</points>
<intersection>365 2</intersection>
<intersection>373 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>365,-199,365,-196.5</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>-199 1</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>371,-195.5,372.5,-195.5</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>363,-202.5,363,-198</points>
<intersection>-202.5 1</intersection>
<intersection>-198 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>363,-202.5,365.5,-202.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>363 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>363,-198,373.5,-198</points>
<intersection>363 0</intersection>
<intersection>373.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>373.5,-198,373.5,-196.5</points>
<connection>
<GID>14</GID>
<name>N_in2</name></connection>
<intersection>-198 2</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>343,-206,347.5,-206</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>340,-193.5,347.5,-193.5</points>
<connection>
<GID>20</GID>
<name>N_in1</name></connection>
<intersection>347.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>347.5,-194,347.5,-193.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-193.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>335,-193.5,338,-193.5</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>20</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>339,-206,339,-194.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-199,347,-196</points>
<connection>
<GID>21</GID>
<name>N_in3</name></connection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>347,-196,347.5,-196</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>347 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,-195,356.5,-194.5</points>
<intersection>-195 2</intersection>
<intersection>-194.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,-194.5,359.5,-194.5</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353.5,-195,356.5,-195</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>356.5,-205,356.5,-204.5</points>
<intersection>-205 2</intersection>
<intersection>-204.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>356.5,-204.5,359.5,-204.5</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>356.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>353.5,-205,356.5,-205</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>356.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>407.5,-196,411,-196</points>
<connection>
<GID>27</GID>
<name>N_in1</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>407.5,-206,411.5,-206</points>
<connection>
<GID>28</GID>
<name>N_in1</name></connection>
<connection>
<GID>26</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>9</ID>
<points>417.5,-205,418,-205</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>29</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>419,-204,419,-200.5</points>
<connection>
<GID>29</GID>
<name>N_in3</name></connection>
<intersection>-200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>411,-200.5,419,-200.5</points>
<intersection>411 2</intersection>
<intersection>419 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>411,-200.5,411,-198</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-200.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>417,-197,418.5,-197</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>409,-204,409,-199.5</points>
<intersection>-204 1</intersection>
<intersection>-199.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>409,-204,411.5,-204</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>409 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>409,-199.5,419.5,-199.5</points>
<intersection>409 0</intersection>
<intersection>419.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>419.5,-199.5,419.5,-198</points>
<connection>
<GID>30</GID>
<name>N_in2</name></connection>
<intersection>-199.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>420.5,-197,424.5,-197</points>
<connection>
<GID>30</GID>
<name>N_in1</name></connection>
<connection>
<GID>31</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>393,-207.5,393.5,-207.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>392,-195.5,393.5,-195.5</points>
<connection>
<GID>42</GID>
<name>N_in1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>389,-207.5,389,-196.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-196.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>389,-196.5,391,-196.5</points>
<connection>
<GID>42</GID>
<name>N_in2</name></connection>
<intersection>389 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,-200.5,393,-197.5</points>
<connection>
<GID>43</GID>
<name>N_in3</name></connection>
<intersection>-197.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>393,-197.5,393.5,-197.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>393 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>393,-205.5,393,-202.5</points>
<connection>
<GID>43</GID>
<name>N_in2</name></connection>
<intersection>-205.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>393,-205.5,393.5,-205.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>393 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-196.5,402.5,-196</points>
<intersection>-196.5 2</intersection>
<intersection>-196 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,-196,405.5,-196</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399.5,-196.5,402.5,-196.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>402.5,-206.5,402.5,-206</points>
<intersection>-206.5 2</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>402.5,-206,405.5,-206</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<intersection>402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399.5,-206.5,402.5,-206.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>347,-216,347,-201</points>
<connection>
<GID>21</GID>
<name>N_in2</name></connection>
<intersection>-216 2</intersection>
<intersection>-204 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>347,-216,361.5,-216</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>347 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>347,-204,347.5,-204</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>347 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>365.5,-216,387,-216</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>370.5 9</intersection>
<intersection>387 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>387,-216,387,-201.5</points>
<intersection>-216 1</intersection>
<intersection>-201.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>387,-201.5,392,-201.5</points>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>387 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>370.5,-220.5,370.5,-216</points>
<connection>
<GID>45</GID>
<name>CLK</name></connection>
<intersection>-216 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>374.5,-195.5,390,-195.5</points>
<connection>
<GID>14</GID>
<name>N_in1</name></connection>
<connection>
<GID>42</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373.5,-194.5,373.5,-191.5</points>
<connection>
<GID>14</GID>
<name>N_in3</name></connection>
<connection>
<GID>46</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>410.5,-242,410.5,-241.5</points>
<intersection>-242 1</intersection>
<intersection>-241.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>409,-242,410.5,-242</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>410.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>410.5,-241.5,412.5,-241.5</points>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<intersection>410.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>401,-242,401,-240.5</points>
<intersection>-242 1</intersection>
<intersection>-240.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>401,-242,403,-242</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>401 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>399,-240.5,401,-240.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>401 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>400.5,-247,400.5,-246</points>
<intersection>-247 2</intersection>
<intersection>-246 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>400.5,-246,403,-246</points>
<connection>
<GID>66</GID>
<name>clock_enable</name></connection>
<intersection>400.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>398,-247,400.5,-247</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>400.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>398,-244,398,-243.5</points>
<intersection>-244 1</intersection>
<intersection>-243.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>398,-244,403,-244</points>
<connection>
<GID>66</GID>
<name>clock</name></connection>
<intersection>398 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>393.5,-243.5,398,-243.5</points>
<connection>
<GID>142</GID>
<name>CLK</name></connection>
<intersection>398 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-86.3,33.2616,51.75,-47.2451</PageViewport>
<gate>
<ID>225</ID>
<type>BB_CLOCK</type>
<position>-56,-39.5</position>
<output>
<ID>CLK</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_TOGGLE</type>
<position>-72,7</position>
<output>
<ID>OUT_0</ID>224 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AA_AND2</type>
<position>-46.5,-13</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AI_XOR2</type>
<position>-46,10</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>254 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>-37.5,5</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>49.5,-3.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>252 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>-21,27</position>
<gparam>LABEL_TEXT 2-bit Counter using D-Latches</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>-20.5,23</position>
<gparam>LABEL_TEXT Should count/output  0,1,2,3,0,..</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>AA_LABEL</type>
<position>18,-7.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>15.5,14.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>AA_LABEL</type>
<position>-73.5,4</position>
<gparam>LABEL_TEXT to enable counter</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>3,-35.5</position>
<gparam>LABEL_TEXT Circuit is not counting correcly</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>-20,-18</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>4,-9</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>BA_NAND2</type>
<position>9.5,-19.5</position>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>6,-21.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>HA_JUNC_2</type>
<position>1.5,-10.5</position>
<input>
<ID>N_in0</ID>235 </input>
<input>
<ID>N_in1</ID>226 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>HA_JUNC_2</type>
<position>1.5,-20.5</position>
<input>
<ID>N_in0</ID>236 </input>
<input>
<ID>N_in1</ID>227 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>HE_JUNC_4</type>
<position>14,-19.5</position>
<input>
<ID>N_in0</ID>228 </input>
<input>
<ID>N_in3</ID>229 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>HE_JUNC_4</type>
<position>14.5,-11.5</position>
<input>
<ID>N_in2</ID>256 </input>
<input>
<ID>N_in3</ID>257 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>-20.5,-10</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>BA_NAND2</type>
<position>-8.5,-11</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>247</ID>
<type>BA_NAND2</type>
<position>-8.5,-21</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AE_SMALL_INVERTER</type>
<position>-14,-22</position>
<input>
<ID>IN_0</ID>232 </input>
<output>
<ID>OUT_0</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>249</ID>
<type>HE_JUNC_4</type>
<position>-14,-10</position>
<input>
<ID>N_in0</ID>237 </input>
<input>
<ID>N_in1</ID>231 </input>
<input>
<ID>N_in2</ID>232 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>BA_NAND2</type>
<position>9.5,-10.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>HE_JUNC_4</type>
<position>-12,-16</position>
<input>
<ID>N_in2</ID>234 </input>
<input>
<ID>N_in3</ID>233 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>-21.5,5</position>
<gparam>LABEL_TEXT WE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AA_LABEL</type>
<position>2.5,14</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>AA_LABEL</type>
<position>4.5,1.5</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>255</ID>
<type>BA_NAND2</type>
<position>7.5,11.5</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>BA_NAND2</type>
<position>8,3.5</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>239 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>HA_JUNC_2</type>
<position>0,12.5</position>
<input>
<ID>N_in0</ID>249 </input>
<input>
<ID>N_in1</ID>238 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>HA_JUNC_2</type>
<position>0,2.5</position>
<input>
<ID>N_in0</ID>250 </input>
<input>
<ID>N_in1</ID>239 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>HE_JUNC_4</type>
<position>12.5,3.5</position>
<input>
<ID>N_in0</ID>240 </input>
<input>
<ID>N_in3</ID>241 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>HE_JUNC_4</type>
<position>13,11.5</position>
<input>
<ID>N_in0</ID>242 </input>
<input>
<ID>N_in1</ID>252 </input>
<input>
<ID>N_in2</ID>243 </input>
<input>
<ID>N_in3</ID>251 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>-22,13</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>BA_NAND2</type>
<position>-10,12</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>BA_NAND2</type>
<position>-10,2</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AE_SMALL_INVERTER</type>
<position>-15.5,1</position>
<input>
<ID>IN_0</ID>246 </input>
<output>
<ID>OUT_0</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>265</ID>
<type>HE_JUNC_4</type>
<position>-15.5,13</position>
<input>
<ID>N_in0</ID>253 </input>
<input>
<ID>N_in1</ID>245 </input>
<input>
<ID>N_in2</ID>246 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>HE_JUNC_4</type>
<position>-13.5,7</position>
<input>
<ID>N_in0</ID>234 </input>
<input>
<ID>N_in2</ID>248 </input>
<input>
<ID>N_in3</ID>247 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AE_SMALL_INVERTER</type>
<position>-52.5,-14</position>
<input>
<ID>IN_0</ID>254 </input>
<output>
<ID>OUT_0</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>-77,10.5</position>
<gparam>LABEL_TEXT "ON" switch</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>274</ID>
<type>AA_LABEL</type>
<position>8.5,-40</position>
<gparam>LABEL_TEXT Problem with using D-latches instead of Flip Flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-59.5,-12,-59.5,7</points>
<intersection>-12 10</intersection>
<intersection>4 12</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-70,7,-59.5,7</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-59.5,-12,-49.5,-12</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-59.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-59.5,4,-40.5,4</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>-59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,6,-42,10</points>
<intersection>6 2</intersection>
<intersection>10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43,10,-42,10</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>-42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,6,-40.5,6</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>-42 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-9.5,6.5,-9.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>2.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>2.5,-10.5,2.5,-9.5</points>
<connection>
<GID>241</GID>
<name>N_in1</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-20.5,6.5,-20.5</points>
<connection>
<GID>242</GID>
<name>N_in1</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-19.5,13,-19.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<connection>
<GID>243</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-18.5,14,-15</points>
<connection>
<GID>243</GID>
<name>N_in3</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,-15,14,-15</points>
<intersection>6 2</intersection>
<intersection>14 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>6,-15,6,-11.5</points>
<intersection>-15 1</intersection>
<intersection>-11.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>6,-11.5,6.5,-11.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>6 2</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-12,-22,-11.5,-22</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,-10,-11.5,-10</points>
<connection>
<GID>249</GID>
<name>N_in1</name></connection>
<connection>
<GID>246</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-22,-16,-11</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16,-11,-14,-11</points>
<connection>
<GID>249</GID>
<name>N_in2</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-15,-12,-12</points>
<connection>
<GID>251</GID>
<name>N_in3</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,-12,-11.5,-12</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,-39.5,-31,7</points>
<intersection>-39.5 5</intersection>
<intersection>-20 1</intersection>
<intersection>-17 6</intersection>
<intersection>7 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31,-20,-11.5,-20</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-31 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-52,-39.5,-31,-39.5</points>
<connection>
<GID>225</GID>
<name>CLK</name></connection>
<intersection>-31 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-31,-17,-12,-17</points>
<connection>
<GID>251</GID>
<name>N_in2</name></connection>
<intersection>-31 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-31,7,-14.5,7</points>
<connection>
<GID>266</GID>
<name>N_in0</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-11,-2.5,-10.5</points>
<intersection>-11 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-10.5,0.5,-10.5</points>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-11,-2.5,-11</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-21,-2.5,-20.5</points>
<intersection>-21 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-20.5,0.5,-20.5</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-21,-2.5,-21</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,-13,-24,-10</points>
<intersection>-13 2</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-10,-15,-10</points>
<connection>
<GID>249</GID>
<name>N_in0</name></connection>
<intersection>-24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43.5,-13,-24,-13</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,12.5,4.5,12.5</points>
<connection>
<GID>257</GID>
<name>N_in1</name></connection>
<connection>
<GID>255</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1,2.5,5,2.5</points>
<connection>
<GID>258</GID>
<name>N_in1</name></connection>
<connection>
<GID>256</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,3.5,11.5,3.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>259</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,4.5,12.5,8</points>
<connection>
<GID>259</GID>
<name>N_in3</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4.5,8,12.5,8</points>
<intersection>4.5 2</intersection>
<intersection>12.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>4.5,8,4.5,10.5</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>8 1</intersection></vsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10.5,11.5,12,11.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<connection>
<GID>260</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,4.5,2.5,9</points>
<intersection>4.5 1</intersection>
<intersection>9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,4.5,5,4.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,9,13,9</points>
<intersection>2.5 0</intersection>
<intersection>13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,9,13,10.5</points>
<connection>
<GID>260</GID>
<name>N_in2</name></connection>
<intersection>9 2</intersection></vsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,1,-13,1</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,13,-13,13</points>
<connection>
<GID>265</GID>
<name>N_in1</name></connection>
<connection>
<GID>262</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,1,-17.5,12</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-17.5,12,-15.5,12</points>
<connection>
<GID>265</GID>
<name>N_in2</name></connection>
<intersection>-17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,8,-13.5,11</points>
<connection>
<GID>266</GID>
<name>N_in3</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,11,-13,11</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,3,-13.5,6</points>
<connection>
<GID>266</GID>
<name>N_in2</name></connection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,3,-13,3</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,12,-4,12.5</points>
<intersection>12 3</intersection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,12.5,-1,12.5</points>
<connection>
<GID>257</GID>
<name>N_in0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7,12,-4,12</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,2,-4,2.5</points>
<intersection>2 3</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,2.5,-1,2.5</points>
<connection>
<GID>258</GID>
<name>N_in0</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7,2,-4,2</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,12.5,13,18</points>
<connection>
<GID>260</GID>
<name>N_in3</name></connection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,18,13,18</points>
<intersection>-49 2</intersection>
<intersection>13 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-49,11,-49,18</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>18 1</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-3.5,30,11.5</points>
<intersection>-3.5 1</intersection>
<intersection>11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-3.5,46.5,-3.5</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,11.5,30,11.5</points>
<connection>
<GID>260</GID>
<name>N_in1</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,5,-25.5,13</points>
<intersection>5 2</intersection>
<intersection>13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,13,-16.5,13</points>
<connection>
<GID>265</GID>
<name>N_in0</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,5,-25.5,5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-31.5,-57.5,9</points>
<intersection>-31.5 2</intersection>
<intersection>-14 5</intersection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,9,-49,9</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57.5,-31.5,21.5,-31.5</points>
<intersection>-57.5 0</intersection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-31.5,21.5,-10.5</points>
<intersection>-31.5 2</intersection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>12.5,-10.5,21.5,-10.5</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<intersection>21.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-57.5,-14,-54.5,-14</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-50.5,-14,-49.5,-14</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-14,14.5,-12.5</points>
<connection>
<GID>244</GID>
<name>N_in2</name></connection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-14,14.5,-14</points>
<intersection>3.5 2</intersection>
<intersection>14.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>3.5,-18.5,3.5,-14</points>
<intersection>-18.5 3</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>3.5,-18.5,6.5,-18.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>3.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-10.5,14.5,-4.5</points>
<connection>
<GID>244</GID>
<name>N_in3</name></connection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-4.5,46.5,-4.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-53.4931,41.7665,51.9931,-19.75</PageViewport>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>13.5,8</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>13.5,22.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AE_DFF_LOW_NT</type>
<position>6.5,17.5</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>151 </output>
<input>
<ID>clock</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_DFF_LOW_NT</type>
<position>6.5,3.5</position>
<input>
<ID>IN_0</ID>149 </input>
<output>
<ID>OUTINV_0</ID>150 </output>
<output>
<ID>OUT_0</ID>148 </output>
<input>
<ID>clock</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>112</ID>
<type>BB_CLOCK</type>
<position>-4,-17.5</position>
<output>
<ID>CLK</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_TOGGLE</type>
<position>-45,21.5</position>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>HA_JUNC_2</type>
<position>-22.5,8.5</position>
<input>
<ID>N_in1</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>23,20</position>
<input>
<ID>N_in0</ID>151 </input>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>23,5.5</position>
<input>
<ID>N_in0</ID>148 </input>
<input>
<ID>N_in1</ID>154 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>-19.5,1.5</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AI_XOR2</type>
<position>-19,24.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_AND2</type>
<position>-10.5,19.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>42.5,13</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>-3,41</position>
<gparam>LABEL_TEXT 2-bit Counter Using Flip Flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-17.5,1.5,16.5</points>
<intersection>-17.5 2</intersection>
<intersection>2.5 1</intersection>
<intersection>16.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,2.5,3.5,2.5</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-17.5,1.5,-17.5</points>
<connection>
<GID>112</GID>
<name>CLK</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>1.5,16.5,3.5,16.5</points>
<connection>
<GID>110</GID>
<name>clock</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,2.5,-32.5,21.5</points>
<intersection>2.5 10</intersection>
<intersection>18.5 12</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-43,21.5,-32.5,21.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-32.5,2.5,-22.5,2.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-32.5,18.5,-13.5,18.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,5.5,10.5,8.5</points>
<intersection>5.5 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,5.5,22,5.5</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,8.5,10.5,8.5</points>
<connection>
<GID>114</GID>
<name>N_in1</name></connection>
<intersection>-22 4</intersection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22,8.5,-22,23.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>8.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,1.5,-6.5,5.5</points>
<intersection>1.5 2</intersection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,5.5,3.5,5.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-16.5,1.5,-6.5,1.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-5,10,2.5</points>
<intersection>-5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22.5,-5,10,-5</points>
<intersection>-22.5 3</intersection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,2.5,10,2.5</points>
<connection>
<GID>111</GID>
<name>OUTINV_0</name></connection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22.5,-5,-22.5,0.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-5 1</intersection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,19.5,10,28.5</points>
<intersection>19.5 1</intersection>
<intersection>20 4</intersection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9.5,19.5,10,19.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-22,28.5,10,28.5</points>
<intersection>-22 3</intersection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22,25.5,-22,28.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>10,20,22,20</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7.5,19.5,3.5,19.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,20.5,-15,24.5</points>
<intersection>20.5 2</intersection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,24.5,-15,24.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>-15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,20.5,-13.5,20.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,5.5,31.5,12</points>
<intersection>5.5 2</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,12,39.5,12</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,5.5,31.5,5.5</points>
<connection>
<GID>116</GID>
<name>N_in1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,13,31.5,20</points>
<intersection>13 2</intersection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,20,31.5,20</points>
<connection>
<GID>115</GID>
<name>N_in1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,13,39.5,13</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-34.4488,51.2665,98.4738,-26.25</PageViewport>
<gate>
<ID>61</ID>
<type>HE_JUNC_4</type>
<position>5.5,-2.5</position>
<input>
<ID>N_in1</ID>53 </input>
<input>
<ID>N_in2</ID>46 </input>
<input>
<ID>N_in3</ID>55 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>HE_JUNC_4</type>
<position>1,43</position>
<input>
<ID>N_in1</ID>30 </input>
<input>
<ID>N_in2</ID>42 </input>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>HE_JUNC_4</type>
<position>1,31</position>
<input>
<ID>N_in0</ID>45 </input>
<input>
<ID>N_in1</ID>43 </input>
<input>
<ID>N_in2</ID>44 </input>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>HE_JUNC_4</type>
<position>4.5,13</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in1</ID>63 </input>
<input>
<ID>N_in2</ID>55 </input>
<input>
<ID>N_in3</ID>68 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>HE_JUNC_4</type>
<position>-1,-14.5</position>
<input>
<ID>N_in0</ID>110 </input>
<input>
<ID>N_in1</ID>69 </input>
<input>
<ID>N_in3</ID>109 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>20.5,50.5</position>
<gparam>LABEL_TEXT Traffic Sign</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>36,42.5</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>36,31</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>15.5,9.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>13.5,-2</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>14.5,-11.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>38,20</position>
<gparam>LABEL_TEXT S0*</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>42,9.5</position>
<gparam>LABEL_TEXT S1*</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>HE_JUNC_4</type>
<position>-3.5,16</position>
<input>
<ID>N_in0</ID>115 </input>
<input>
<ID>N_in1</ID>112 </input>
<input>
<ID>N_in2</ID>110 </input>
<input>
<ID>N_in3</ID>113 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>HA_JUNC_2</type>
<position>-3,38.5</position>
<input>
<ID>N_in0</ID>115 </input>
<input>
<ID>N_in1</ID>114 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>HE_JUNC_4</type>
<position>20.5,30.5</position>
<input>
<ID>N_in0</ID>121 </input>
<input>
<ID>N_in2</ID>123 </input>
<input>
<ID>N_in3</ID>122 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>HE_JUNC_4</type>
<position>26,29.5</position>
<input>
<ID>N_in0</ID>137 </input>
<input>
<ID>N_in1</ID>126 </input>
<input>
<ID>N_in2</ID>125 </input>
<input>
<ID>N_in3</ID>127 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>HE_JUNC_4</type>
<position>23.5,27.5</position>
<input>
<ID>N_in1</ID>129 </input>
<input>
<ID>N_in2</ID>130 </input>
<input>
<ID>N_in3</ID>128 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>HE_JUNC_4</type>
<position>24,16</position>
<input>
<ID>N_in0</ID>131 </input>
<input>
<ID>N_in1</ID>132 </input>
<input>
<ID>N_in2</ID>133 </input>
<input>
<ID>N_in3</ID>130 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>HE_JUNC_4</type>
<position>53.5,40</position>
<input>
<ID>N_in0</ID>136 </input>
<input>
<ID>N_in1</ID>134 </input>
<input>
<ID>N_in2</ID>135 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>HE_JUNC_4</type>
<position>65,16.5</position>
<input>
<ID>N_in0</ID>138 </input>
<input>
<ID>N_in1</ID>140 </input>
<input>
<ID>N_in3</ID>139 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>BB_CLOCK</type>
<position>17.5,-24</position>
<output>
<ID>CLK</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>88</ID>
<type>HE_JUNC_4</type>
<position>25.5,-24</position>
<input>
<ID>N_in0</ID>141 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>HE_JUNC_4</type>
<position>25.5,-17</position>
<input>
<ID>N_in0</ID>142 </input>
<input>
<ID>N_in2</ID>141 </input>
<input>
<ID>N_in3</ID>143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>56,31.5</position>
<input>
<ID>N_in3</ID>134 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>GA_LED</type>
<position>56,21</position>
<input>
<ID>N_in3</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>65,28</position>
<input>
<ID>N_in1</ID>140 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>65,23.5</position>
<input>
<ID>N_in2</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>74.5,25.5</position>
<input>
<ID>N_in2</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND3</type>
<position>11.5,40.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>27 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND3</type>
<position>12,29</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>113 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND3</type>
<position>11.5,18</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>63 </input>
<input>
<ID>IN_2</ID>29 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_AND3</type>
<position>11.5,7.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>53 </input>
<input>
<ID>IN_2</ID>109 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_OR3</type>
<position>32,40</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>128 </input>
<input>
<ID>IN_2</ID>127 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_OR2</type>
<position>32,28.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_OR2</type>
<position>32.5,17</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_OR2</type>
<position>33,7.5</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>5.5,40.5</position>
<input>
<ID>IN_0</ID>120 </input>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>5.5,38.5</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_SMALL_INVERTER</type>
<position>6.5,29</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_SMALL_INVERTER</type>
<position>0,16</position>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_DFF_LOW</type>
<position>20,-3</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_DFF_LOW</type>
<position>20,-12.5</position>
<input>
<ID>IN_0</ID>145 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>142 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>-10.5,43</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,40.5,8.5,40.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7.5,38.5,8.5,38.5</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,29,9,29</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<connection>
<GID>96</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,16,8.5,16</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>97</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,42.5,5,43</points>
<intersection>42.5 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5,42.5,8.5,42.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,43,5,43</points>
<connection>
<GID>62</GID>
<name>N_in1</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,43,1,44</points>
<connection>
<GID>62</GID>
<name>N_in3</name></connection>
<intersection>43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,43,1,43</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,32,1,42</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<connection>
<GID>62</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>2,31,9,31</points>
<connection>
<GID>68</GID>
<name>N_in1</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,20,1,30</points>
<connection>
<GID>68</GID>
<name>N_in2</name></connection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,20,8.5,20</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,9.5,2.5,31</points>
<intersection>9.5 1</intersection>
<intersection>31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,9.5,8.5,9.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,31,2.5,31</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-5,5.5,-3.5</points>
<connection>
<GID>61</GID>
<name>N_in2</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-5,17,-5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-2.5,7.5,7.5</points>
<intersection>-2.5 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,7.5,8.5,7.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-2.5,7.5,-2.5</points>
<connection>
<GID>61</GID>
<name>N_in1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-1.5,4.5,12</points>
<connection>
<GID>69</GID>
<name>N_in2</name></connection>
<intersection>-1.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>4.5,-1.5,5.5,-1.5</points>
<connection>
<GID>61</GID>
<name>N_in3</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,13,7.5,18</points>
<intersection>13 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,18,8.5,18</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5.5,13,7.5,13</points>
<connection>
<GID>69</GID>
<name>N_in1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,14,4.5,29</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-14.5,17,-14.5</points>
<connection>
<GID>70</GID>
<name>N_in1</name></connection>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-13.5,-1,5.5</points>
<connection>
<GID>70</GID>
<name>N_in3</name></connection>
<intersection>5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,5.5,8.5,5.5</points>
<connection>
<GID>98</GID>
<name>IN_2</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-14.5,-3.5,15</points>
<connection>
<GID>79</GID>
<name>N_in2</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-14.5,-2,-14.5</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-2.5,16,-2,16</points>
<connection>
<GID>79</GID>
<name>N_in1</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,17,-3.5,27</points>
<connection>
<GID>79</GID>
<name>N_in3</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,27,9,27</points>
<connection>
<GID>96</GID>
<name>IN_2</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-2,38.5,3.5,38.5</points>
<connection>
<GID>80</GID>
<name>N_in1</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,16,-4.5,38.5</points>
<connection>
<GID>79</GID>
<name>N_in0</name></connection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,38.5,-4,38.5</points>
<connection>
<GID>80</GID>
<name>N_in0</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,13,3.5,40.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,29,17,30.5</points>
<intersection>29 2</intersection>
<intersection>30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,30.5,19.5,30.5</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,29,17,29</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,31.5,20.5,42</points>
<connection>
<GID>81</GID>
<name>N_in3</name></connection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,42,29,42</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,18,20.5,29.5</points>
<connection>
<GID>81</GID>
<name>N_in2</name></connection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,18,29.5,18</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,6.5,17.5,40.5</points>
<intersection>6.5 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,40.5,17.5,40.5</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,6.5,30,6.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,7.5,26,28.5</points>
<connection>
<GID>82</GID>
<name>N_in2</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,7.5,26,7.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>27,29.5,29,29.5</points>
<connection>
<GID>82</GID>
<name>N_in1</name></connection>
<connection>
<GID>100</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,30.5,26,38</points>
<connection>
<GID>82</GID>
<name>N_in3</name></connection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,38,29,38</points>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,28.5,23.5,40</points>
<connection>
<GID>83</GID>
<name>N_in3</name></connection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,40,29,40</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>24.5,27.5,29,27.5</points>
<connection>
<GID>83</GID>
<name>N_in1</name></connection>
<connection>
<GID>100</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,22,23.5,26.5</points>
<connection>
<GID>83</GID>
<name>N_in2</name></connection>
<intersection>22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>24,17,24,22</points>
<connection>
<GID>84</GID>
<name>N_in3</name></connection>
<intersection>22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,22,24,22</points>
<intersection>23.5 0</intersection>
<intersection>24 1</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,16,18.5,18</points>
<intersection>16 2</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,18,18.5,18</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,16,23,16</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>25,16,29.5,16</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<connection>
<GID>101</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,8.5,24,15</points>
<connection>
<GID>84</GID>
<name>N_in2</name></connection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,8.5,30,8.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,32.5,56,40</points>
<connection>
<GID>90</GID>
<name>N_in3</name></connection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,40,56,40</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,22,53.5,39</points>
<connection>
<GID>85</GID>
<name>N_in2</name></connection>
<intersection>22 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>53.5,22,56,22</points>
<connection>
<GID>91</GID>
<name>N_in3</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,40,52.5,40</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,24.5,74.5,35</points>
<connection>
<GID>94</GID>
<name>N_in2</name></connection>
<intersection>35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,35,74.5,35</points>
<intersection>25 2</intersection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>25,29.5,25,35</points>
<connection>
<GID>82</GID>
<name>N_in0</name></connection>
<intersection>35 1</intersection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,16.5,49.5,28.5</points>
<intersection>16.5 1</intersection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,16.5,64,16.5</points>
<connection>
<GID>86</GID>
<name>N_in0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,28.5,49.5,28.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,17.5,65,22.5</points>
<connection>
<GID>86</GID>
<name>N_in3</name></connection>
<connection>
<GID>93</GID>
<name>N_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,16.5,67,28</points>
<intersection>16.5 2</intersection>
<intersection>28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,28,67,28</points>
<connection>
<GID>92</GID>
<name>N_in1</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66,16.5,67,16.5</points>
<connection>
<GID>86</GID>
<name>N_in1</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>21.5,-24,25.5,-24</points>
<connection>
<GID>87</GID>
<name>CLK</name></connection>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>25.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>25.5,-24,25.5,-18</points>
<connection>
<GID>89</GID>
<name>N_in2</name></connection>
<intersection>-24 5</intersection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-17,23.5,-11.5</points>
<intersection>-17 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-11.5,23.5,-11.5</points>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-17,24.5,-17</points>
<connection>
<GID>89</GID>
<name>N_in0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-16,25.5,-2</points>
<connection>
<GID>89</GID>
<name>N_in3</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-2,25.5,-2</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-5,38.5,17</points>
<intersection>-5 2</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,17,38.5,17</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-5,38.5,-5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-14.5,42.5,7.5</points>
<intersection>-14.5 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,7.5,42.5,7.5</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-14.5,42.5,-14.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-0.428691,0.25,8.08798,-4.71667</PageViewport></page 4>
<page 5>
<PageViewport>-1e+010,-117.734,-1e+010,-187.25</PageViewport></page 5>
<page 6>
<PageViewport>-1e+010,35.5588,-1e+010,-560.441</PageViewport></page 6>
<page 7>
<PageViewport>-882.076,1283.77,139.924,687.767</PageViewport></page 7>
<page 8>
<PageViewport>-1e+010,-73.233,-1e+010,-669.233</PageViewport></page 8>
<page 9>
<PageViewport>-1e+010,-314.725,-1e+010,-432.167</PageViewport></page 9></circuit>