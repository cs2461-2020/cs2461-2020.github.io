<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-87.9116,54.7665,-6.2131,5.48381</PageViewport>
<gate>
<ID>193</ID>
<type>VE_PMOS</type>
<position>-64.5,42.5</position>
<input>
<ID>T_ctrl</ID>87 </input>
<input>
<ID>T_in</ID>88 </input>
<input>
<ID>T_in2</ID>82 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>194</ID>
<type>VE_PMOS</type>
<position>-57.5,43</position>
<input>
<ID>T_ctrl</ID>86 </input>
<input>
<ID>T_in</ID>88 </input>
<input>
<ID>T_in2</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>2</ID>
<type>VE_PMOS</type>
<position>-28,21</position>
<input>
<ID>T_ctrl</ID>3 </input>
<input>
<ID>T_in</ID>13 </input>
<input>
<ID>T_in2</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>195</ID>
<type>VA_NMOS</type>
<position>-64.5,34</position>
<input>
<ID>T_ctrl</ID>86 </input>
<input>
<ID>T_in</ID>84 </input>
<input>
<ID>T_in2</ID>88 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>-59,54</position>
<gparam>LABEL_TEXT NAND Gate and NOT Gates</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>-43.5,48</position>
<gparam>LABEL_TEXT Parallel circuit on top</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>-47.5,35</position>
<gparam>LABEL_TEXT Series circuit on bottom</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>VA_NMOS</type>
<position>-83,18.5</position>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>10</ID>
<type>VA_NMOS</type>
<position>-28,16</position>
<input>
<ID>T_ctrl</ID>3 </input>
<input>
<ID>T_in</ID>11 </input>
<input>
<ID>T_in2</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>203</ID>
<type>VE_PMOS</type>
<position>-64,17.5</position>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>11</ID>
<type>EE_VDD</type>
<position>-27,26.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>-23.5,28.5</position>
<gparam>LABEL_TEXT Power: 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>FF_GND</type>
<position>-27,12</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>-17,18.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>-15.5,15.5</position>
<gparam>LABEL_TEXT Output Y = NOT X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>-81,21</position>
<gparam>LABEL_TEXT N-type Transistor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>-62.5,21</position>
<gparam>LABEL_TEXT P-type Transistor</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-45.5,18</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-45,20.5</position>
<gparam>LABEL_TEXT Input X</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>VA_NMOS</type>
<position>-64.5,30.5</position>
<input>
<ID>T_ctrl</ID>87 </input>
<input>
<ID>T_in</ID>83 </input>
<input>
<ID>T_in2</ID>84 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_TOGGLE</type>
<position>-72.5,42.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>-72.5,38.5</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>-75,43</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>-76,38.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>181</ID>
<type>GA_LED</type>
<position>-52,38.5</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>-52.5,41.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>183</ID>
<type>EE_VDD</type>
<position>-63.5,47.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-54.5,50</position>
<gparam>LABEL_TEXT Power: 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>FF_GND</type>
<position>-63.5,26.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-59,27</position>
<gparam>LABEL_TEXT Ground: 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>EE_VDD</type>
<position>-56.5,47.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>-42.5,46</position>
<gparam>LABEL_TEXT If one of the top two closes</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>-40.5,44.5</position>
<gparam>LABEL_TEXT then connection to power and C=1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>-48.5,33</position>
<gparam>LABEL_TEXT If both lower two transistors close</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>-48,31.5</position>
<gparam>LABEL_TEXT then connection to ground and C=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>-39,16,-39,21</points>
<intersection>16 12</intersection>
<intersection>18 13</intersection>
<intersection>21 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-39,21,-30,21</points>
<connection>
<GID>2</GID>
<name>T_ctrl</name></connection>
<intersection>-39 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-39,16,-30,16</points>
<connection>
<GID>10</GID>
<name>T_ctrl</name></connection>
<intersection>-39 9</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-43.5,18,-39,18</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-39 9</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,13,-27,15</points>
<connection>
<GID>10</GID>
<name>T_in</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,22,-27,25.5</points>
<connection>
<GID>2</GID>
<name>T_in2</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,17,-27,20</points>
<connection>
<GID>10</GID>
<name>T_in2</name></connection>
<connection>
<GID>2</GID>
<name>T_in</name></connection>
<intersection>18.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-27,18.5,-18,18.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,43.5,-63.5,46.5</points>
<connection>
<GID>193</GID>
<name>T_in2</name></connection>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,27.5,-63.5,29.5</points>
<connection>
<GID>176</GID>
<name>T_in</name></connection>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,31.5,-63.5,33</points>
<connection>
<GID>176</GID>
<name>T_in2</name></connection>
<connection>
<GID>195</GID>
<name>T_in</name></connection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,44,-56.5,46.5</points>
<connection>
<GID>194</GID>
<name>T_in2</name></connection>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,34,-68.5,49</points>
<intersection>34 1</intersection>
<intersection>42.5 2</intersection>
<intersection>49 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,34,-66.5,34</points>
<connection>
<GID>195</GID>
<name>T_ctrl</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,42.5,-68.5,42.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-68.5,49,-59.5,49</points>
<intersection>-68.5 0</intersection>
<intersection>-59.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-59.5,43,-59.5,49</points>
<connection>
<GID>194</GID>
<name>T_ctrl</name></connection>
<intersection>49 3</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69.5,30.5,-69.5,40.5</points>
<intersection>30.5 1</intersection>
<intersection>38.5 2</intersection>
<intersection>40.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69.5,30.5,-66.5,30.5</points>
<connection>
<GID>176</GID>
<name>T_ctrl</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-70.5,38.5,-69.5,38.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>-69.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-69.5,40.5,-66.5,40.5</points>
<intersection>-69.5 0</intersection>
<intersection>-66.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-66.5,40.5,-66.5,42.5</points>
<connection>
<GID>193</GID>
<name>T_ctrl</name></connection>
<intersection>40.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60,35,-60,38.5</points>
<intersection>35 4</intersection>
<intersection>38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-63.5,38.5,-53,38.5</points>
<connection>
<GID>181</GID>
<name>N_in0</name></connection>
<intersection>-63.5 7</intersection>
<intersection>-60 0</intersection>
<intersection>-56.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-63.5,35,-60,35</points>
<connection>
<GID>195</GID>
<name>T_in2</name></connection>
<intersection>-60 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-56.5,38.5,-56.5,42</points>
<connection>
<GID>194</GID>
<name>T_in</name></connection>
<intersection>38.5 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-63.5,38.5,-63.5,41.5</points>
<connection>
<GID>193</GID>
<name>T_in</name></connection>
<intersection>38.5 3</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-21.2957,52.5082,37.7695,16.8785</PageViewport>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>-3.5,52</position>
<gparam>LABEL_TEXT Question</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>AA_LABEL</type>
<position>-4.5,50</position>
<gparam>LABEL_TEXT Which gate is being  implemented ?</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_LABEL</type>
<position>15,29</position>
<gparam>LABEL_TEXT If one of the bottom two closes</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_LABEL</type>
<position>17,27.5</position>
<gparam>LABEL_TEXT then connection to ground and C=0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>10.5,41</position>
<gparam>LABEL_TEXT If both upper two transistors close</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>11,39.5</position>
<gparam>LABEL_TEXT then connection to power and C=1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>VE_PMOS</type>
<position>-5,40.5</position>
<input>
<ID>T_ctrl</ID>79 </input>
<input>
<ID>T_in</ID>76 </input>
<input>
<ID>T_in2</ID>80 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>162</ID>
<type>VE_PMOS</type>
<position>-5,35.5</position>
<input>
<ID>T_ctrl</ID>78 </input>
<input>
<ID>T_in</ID>77 </input>
<input>
<ID>T_in2</ID>76 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>163</ID>
<type>VA_NMOS</type>
<position>-7,28.5</position>
<input>
<ID>T_ctrl</ID>79 </input>
<input>
<ID>T_in</ID>81 </input>
<input>
<ID>T_in2</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>164</ID>
<type>VA_NMOS</type>
<position>0.5,28.5</position>
<input>
<ID>T_ctrl</ID>78 </input>
<input>
<ID>T_in</ID>81 </input>
<input>
<ID>T_in2</ID>77 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_TOGGLE</type>
<position>-13.5,40.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>-13.5,35.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>-15.5,41</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>-15.5,36</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>6.5,33.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>6,35.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>171</ID>
<type>EE_VDD</type>
<position>-4,45</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>0,47</position>
<gparam>LABEL_TEXT Power: 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>FF_GND</type>
<position>-4,22.5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>0.5,22</position>
<gparam>LABEL_TEXT Ground: 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,36.5,-4,39.5</points>
<connection>
<GID>162</GID>
<name>T_in2</name></connection>
<connection>
<GID>161</GID>
<name>T_in</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,32,2,32</points>
<intersection>-6 6</intersection>
<intersection>-4 3</intersection>
<intersection>2 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-4,32,-4,34.5</points>
<connection>
<GID>162</GID>
<name>T_in</name></connection>
<intersection>32 1</intersection>
<intersection>33.5 10</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>2,29.5,2,32</points>
<intersection>29.5 8</intersection>
<intersection>32 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-6,29.5,-6,32</points>
<connection>
<GID>163</GID>
<name>T_in2</name></connection>
<intersection>32 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>1.5,29.5,2,29.5</points>
<connection>
<GID>164</GID>
<name>T_in2</name></connection>
<intersection>2 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-4,33.5,5.5,33.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<intersection>-4 3</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,35.5,-7,35.5</points>
<connection>
<GID>162</GID>
<name>T_ctrl</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,25,-11.5,35.5</points>
<intersection>25 4</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11.5,25,-3,25</points>
<intersection>-11.5 3</intersection>
<intersection>-3 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-3,25,-3,28.5</points>
<intersection>25 4</intersection>
<intersection>28.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-3,28.5,-1.5,28.5</points>
<connection>
<GID>164</GID>
<name>T_ctrl</name></connection>
<intersection>-3 5</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,40.5,-7,40.5</points>
<connection>
<GID>161</GID>
<name>T_ctrl</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,28.5,-11.5,40.5</points>
<intersection>28.5 5</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-11.5,28.5,-9,28.5</points>
<connection>
<GID>163</GID>
<name>T_ctrl</name></connection>
<intersection>-11.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,41.5,-4,44</points>
<connection>
<GID>161</GID>
<name>T_in2</name></connection>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,23.5,1.5,23.5</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>-6 3</intersection>
<intersection>1.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>1.5,23.5,1.5,27.5</points>
<connection>
<GID>164</GID>
<name>T_in</name></connection>
<intersection>23.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>-6,23.5,-6,27.5</points>
<connection>
<GID>163</GID>
<name>T_in</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>113.424,-40.9918,171.501,-76.025</PageViewport>
<gate>
<ID>1</ID>
<type>VE_PMOS</type>
<position>127.5,-56.5</position>
<input>
<ID>T_ctrl</ID>7 </input>
<input>
<ID>T_in</ID>4 </input>
<input>
<ID>T_in2</ID>8 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>3</ID>
<type>VE_PMOS</type>
<position>127.5,-61.5</position>
<input>
<ID>T_ctrl</ID>6 </input>
<input>
<ID>T_in</ID>5 </input>
<input>
<ID>T_in2</ID>4 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>4</ID>
<type>VA_NMOS</type>
<position>125.5,-68.5</position>
<input>
<ID>T_ctrl</ID>7 </input>
<input>
<ID>T_in</ID>9 </input>
<input>
<ID>T_in2</ID>5 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>5</ID>
<type>VA_NMOS</type>
<position>133,-68.5</position>
<input>
<ID>T_ctrl</ID>6 </input>
<input>
<ID>T_in</ID>9 </input>
<input>
<ID>T_in2</ID>5 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>119,-56.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>119,-61.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>117,-56</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>117,-61</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>12</ID>
<type>EE_VDD</type>
<position>128.5,-52</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>13</ID>
<type>FF_GND</type>
<position>128.5,-74.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>133,-75</position>
<gparam>LABEL_TEXT Ground: 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>VE_PMOS</type>
<position>152.5,-61</position>
<input>
<ID>T_ctrl</ID>10 </input>
<input>
<ID>T_in</ID>55 </input>
<input>
<ID>T_in2</ID>54 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>16</ID>
<type>VA_NMOS</type>
<position>152.5,-66</position>
<input>
<ID>T_ctrl</ID>10 </input>
<input>
<ID>T_in</ID>53 </input>
<input>
<ID>T_in2</ID>55 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>17</ID>
<type>EE_VDD</type>
<position>153.5,-55.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>FF_GND</type>
<position>153.5,-70</position>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>163.5,-63.5</position>
<input>
<ID>N_in0</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>165,-66.5</position>
<gparam>LABEL_TEXT Output D</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>HA_JUNC_2</type>
<position>135,-63</position>
<input>
<ID>N_in0</ID>5 </input>
<input>
<ID>N_in1</ID>10 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>141.5,-44</position>
<gparam>LABEL_TEXT Combining gates to build new 'gates'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>129,-50</position>
<gparam>LABEL_TEXT This part is gate from page 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>142,-41.5</position>
<gparam>LABEL_TEXT Which gate is being  implemented ?</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-60.5,128.5,-57.5</points>
<connection>
<GID>3</GID>
<name>T_in2</name></connection>
<connection>
<GID>1</GID>
<name>T_in</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126.5,-65,134.5,-65</points>
<intersection>126.5 6</intersection>
<intersection>128.5 3</intersection>
<intersection>134.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-65,128.5,-62.5</points>
<connection>
<GID>3</GID>
<name>T_in</name></connection>
<intersection>-65 1</intersection>
<intersection>-63 14</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>134.5,-67.5,134.5,-65</points>
<intersection>-67.5 8</intersection>
<intersection>-65 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>126.5,-67.5,126.5,-65</points>
<connection>
<GID>4</GID>
<name>T_in2</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>134,-67.5,134.5,-67.5</points>
<connection>
<GID>5</GID>
<name>T_in2</name></connection>
<intersection>134.5 5</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>128.5,-63,134,-63</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>128.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121,-61.5,125.5,-61.5</points>
<connection>
<GID>3</GID>
<name>T_ctrl</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121,-72,121,-61.5</points>
<intersection>-72 4</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>121,-72,129.5,-72</points>
<intersection>121 3</intersection>
<intersection>129.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>129.5,-72,129.5,-68.5</points>
<intersection>-72 4</intersection>
<intersection>-68.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>129.5,-68.5,131,-68.5</points>
<connection>
<GID>5</GID>
<name>T_ctrl</name></connection>
<intersection>129.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121,-56.5,125.5,-56.5</points>
<connection>
<GID>1</GID>
<name>T_ctrl</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>121 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121,-68.5,121,-56.5</points>
<intersection>-68.5 5</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>121,-68.5,123.5,-68.5</points>
<connection>
<GID>4</GID>
<name>T_ctrl</name></connection>
<intersection>121 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128.5,-55.5,128.5,-53</points>
<connection>
<GID>1</GID>
<name>T_in2</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>126.5,-73.5,134,-73.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>126.5 3</intersection>
<intersection>134 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>134,-73.5,134,-69.5</points>
<connection>
<GID>5</GID>
<name>T_in</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>126.5,-73.5,126.5,-69.5</points>
<connection>
<GID>4</GID>
<name>T_in</name></connection>
<intersection>-73.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>141.5,-66,141.5,-61</points>
<intersection>-66 12</intersection>
<intersection>-63 13</intersection>
<intersection>-61 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>141.5,-61,150.5,-61</points>
<connection>
<GID>15</GID>
<name>T_ctrl</name></connection>
<intersection>141.5 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>141.5,-66,150.5,-66</points>
<connection>
<GID>16</GID>
<name>T_ctrl</name></connection>
<intersection>141.5 9</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>136,-63,141.5,-63</points>
<connection>
<GID>22</GID>
<name>N_in1</name></connection>
<intersection>141.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-69,153.5,-67</points>
<connection>
<GID>16</GID>
<name>T_in</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-60,153.5,-56.5</points>
<connection>
<GID>15</GID>
<name>T_in2</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-65,153.5,-62</points>
<connection>
<GID>16</GID>
<name>T_in2</name></connection>
<connection>
<GID>15</GID>
<name>T_in</name></connection>
<intersection>-63.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>153.5,-63.5,162.5,-63.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>39.296,177.953,141.229,116.464</PageViewport>
<gate>
<ID>34</ID>
<type>VE_PMOS</type>
<position>78,156.5</position>
<input>
<ID>T_ctrl</ID>14 </input>
<input>
<ID>T_in</ID>17 </input>
<input>
<ID>T_in2</ID>16 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>35</ID>
<type>VA_NMOS</type>
<position>78,151.5</position>
<input>
<ID>T_ctrl</ID>14 </input>
<input>
<ID>T_in</ID>15 </input>
<input>
<ID>T_in2</ID>17 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>36</ID>
<type>EE_VDD</type>
<position>79,162</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>37</ID>
<type>FF_GND</type>
<position>79,147.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>82.5,156</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>VE_PMOS</type>
<position>78,134.5</position>
<input>
<ID>T_ctrl</ID>18 </input>
<input>
<ID>T_in</ID>21 </input>
<input>
<ID>T_in2</ID>20 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>55</ID>
<type>VA_NMOS</type>
<position>78,129.5</position>
<input>
<ID>T_ctrl</ID>18 </input>
<input>
<ID>T_in</ID>19 </input>
<input>
<ID>T_in2</ID>21 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>59</ID>
<type>EE_VDD</type>
<position>79,140</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>FF_GND</type>
<position>79,125.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>82.5,130.5</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>84,169.5</position>
<gparam>LABEL_TEXT Find Truth Table for C,D,F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>62.5,154.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>63.5,132.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>VE_PMOS</type>
<position>98,154</position>
<input>
<ID>T_ctrl</ID>65 </input>
<input>
<ID>T_in</ID>56 </input>
<input>
<ID>T_in2</ID>60 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>66,154</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>67,132</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>114</ID>
<type>VE_PMOS</type>
<position>98,149</position>
<input>
<ID>T_ctrl</ID>66 </input>
<input>
<ID>T_in</ID>67 </input>
<input>
<ID>T_in2</ID>56 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>115</ID>
<type>VA_NMOS</type>
<position>93.5,139.5</position>
<input>
<ID>T_ctrl</ID>65 </input>
<input>
<ID>T_in</ID>63 </input>
<input>
<ID>T_in2</ID>67 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>116</ID>
<type>VA_NMOS</type>
<position>98,132</position>
<input>
<ID>T_ctrl</ID>66 </input>
<input>
<ID>T_in</ID>62 </input>
<input>
<ID>T_in2</ID>67 </input>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>121</ID>
<type>EE_VDD</type>
<position>99,162.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>122</ID>
<type>FF_GND</type>
<position>102.5,126.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>HA_JUNC_2</type>
<position>105.5,144</position>
<input>
<ID>N_in0</ID>67 </input>
<input>
<ID>N_in1</ID>68 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>82.5,154</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>82.5,132</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>74.5,166.5</position>
<gparam>LABEL_TEXT Ground: 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>FF_GND</type>
<position>79.5,166</position>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>EE_VDD</type>
<position>92.5,166.5</position>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>87.5,166.5</position>
<gparam>LABEL_TEXT Power: 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>FF_GND</type>
<position>94.5,135.5</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>109.5,144</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>112,145</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>72,151.5,72,156.5</points>
<intersection>151.5 12</intersection>
<intersection>154 13</intersection>
<intersection>156.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>72,156.5,76,156.5</points>
<connection>
<GID>34</GID>
<name>T_ctrl</name></connection>
<intersection>72 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>72,151.5,76,151.5</points>
<connection>
<GID>35</GID>
<name>T_ctrl</name></connection>
<intersection>72 9</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>68,154,72,154</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>72 9</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,148.5,79,150.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<connection>
<GID>35</GID>
<name>T_in</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,157.5,79,161</points>
<connection>
<GID>34</GID>
<name>T_in2</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,152.5,79,155.5</points>
<connection>
<GID>35</GID>
<name>T_in2</name></connection>
<connection>
<GID>34</GID>
<name>T_in</name></connection>
<intersection>154 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>79,154,81.5,154</points>
<connection>
<GID>127</GID>
<name>N_in0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>9</ID>
<points>72,129.5,72,134.5</points>
<intersection>129.5 12</intersection>
<intersection>132 13</intersection>
<intersection>134.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>72,134.5,76,134.5</points>
<connection>
<GID>53</GID>
<name>T_ctrl</name></connection>
<intersection>72 9</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>72,129.5,76,129.5</points>
<connection>
<GID>55</GID>
<name>T_ctrl</name></connection>
<intersection>72 9</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>69,132,72,132</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>72 9</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,126.5,79,128.5</points>
<connection>
<GID>55</GID>
<name>T_in</name></connection>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,135.5,79,139</points>
<connection>
<GID>53</GID>
<name>T_in2</name></connection>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,130.5,79,133.5</points>
<connection>
<GID>53</GID>
<name>T_in</name></connection>
<connection>
<GID>55</GID>
<name>T_in2</name></connection>
<intersection>132 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>79,132,81.5,132</points>
<connection>
<GID>129</GID>
<name>N_in0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,150,99,153</points>
<connection>
<GID>114</GID>
<name>T_in2</name></connection>
<connection>
<GID>103</GID>
<name>T_in</name></connection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>99,155,99,161.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<connection>
<GID>103</GID>
<name>T_in2</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,127.5,99,131</points>
<connection>
<GID>116</GID>
<name>T_in</name></connection>
<intersection>127.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>99,127.5,102.5,127.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,136.5,94.5,138.5</points>
<connection>
<GID>115</GID>
<name>T_in</name></connection>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83.5,154,96,154</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<connection>
<GID>103</GID>
<name>T_ctrl</name></connection>
<intersection>90 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>90,139.5,90,154</points>
<intersection>139.5 5</intersection>
<intersection>154 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>90,139.5,91.5,139.5</points>
<connection>
<GID>115</GID>
<name>T_ctrl</name></connection>
<intersection>90 4</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,132,96,132</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<connection>
<GID>116</GID>
<name>T_ctrl</name></connection>
<intersection>82.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>82.5,132,82.5,149</points>
<intersection>132 1</intersection>
<intersection>149 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>82.5,149,96,149</points>
<connection>
<GID>114</GID>
<name>T_ctrl</name></connection>
<intersection>82.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,133,99,148</points>
<connection>
<GID>116</GID>
<name>T_in2</name></connection>
<connection>
<GID>114</GID>
<name>T_in</name></connection>
<intersection>144 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>94.5,144,104.5,144</points>
<connection>
<GID>124</GID>
<name>N_in0</name></connection>
<intersection>94.5 5</intersection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>94.5,140.5,94.5,144</points>
<connection>
<GID>115</GID>
<name>T_in2</name></connection>
<intersection>144 4</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>106.5,144,108.5,144</points>
<connection>
<GID>124</GID>
<name>N_in1</name></connection>
<connection>
<GID>138</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-87.25,58.6181,-17.4396,16.5067</PageViewport>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>-48.5,43</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>-48.5,40</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_OR2</type>
<position>-39,32</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_TOGGLE</type>
<position>-48,30</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-86,43.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-86,40.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-85.5,32.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-85.5,29</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-52,43.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>-52,40.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-52,30.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-41,48.5</position>
<gparam>LABEL_TEXT (A AND B) AND ( NOT B OR C)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>-73,41.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>-81.5,43</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>-81.5,40</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>-64,41.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AE_OR2</type>
<position>-72,30.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_TOGGLE</type>
<position>-81,31.5</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>-81,28.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>106</ID>
<type>GA_LED</type>
<position>-62.5,30.5</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AE_SMALL_INVERTER</type>
<position>-44,33</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>-30.5,37.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>-23.5,37.5</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>-76.5,52</position>
<gparam>LABEL_TEXT Examples</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>-75,46.5</position>
<gparam>LABEL_TEXT A AND B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>-74.5,35</position>
<gparam>LABEL_TEXT A OR B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>-40,41.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-42,33,-42,33</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,38.5,-35,41.5</points>
<intersection>38.5 1</intersection>
<intersection>41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,38.5,-33.5,38.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37,41.5,-35,41.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34.5,32,-34.5,36.5</points>
<intersection>32 1</intersection>
<intersection>36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,32,-34.5,32</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-34.5,36.5,-33.5,36.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,37.5,-24.5,37.5</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,42.5,-44.5,43</points>
<intersection>42.5 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,42.5,-43,42.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46.5,43,-44.5,43</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,40,-44.5,40.5</points>
<intersection>40 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,40.5,-43,40.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46.5,40,-44.5,40</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 3</intersection>
<intersection>-44.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-46.5,33,-46.5,40</points>
<intersection>33 4</intersection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-46.5,33,-46,33</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-46.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,30,-44,31</points>
<intersection>30 2</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44,31,-42,31</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46,30,-44,30</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-70,41.5,-65,41.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,42.5,-77.5,43</points>
<intersection>42.5 1</intersection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,42.5,-76,42.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,43,-77.5,43</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,40,-77.5,40.5</points>
<intersection>40 2</intersection>
<intersection>40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,40.5,-76,40.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,40,-77.5,40</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-79,31.5,-75,31.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77,28.5,-77,29.5</points>
<intersection>28.5 2</intersection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77,29.5,-75,29.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>-77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79,28.5,-77,28.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-77 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-69,30.5,-63.5,30.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>392.277,37.7665,479.502,-14.8494</PageViewport>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>438,6.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>433,37</position>
<gparam>LABEL_TEXT (a) What is the boolean function for this circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>433,32.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>415.5,33.5</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>47</ID>
<type>AE_SMALL_INVERTER</type>
<position>424.5,31.5</position>
<input>
<ID>IN_0</ID>32 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>433.5,23.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_SMALL_INVERTER</type>
<position>426.5,24.5</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>415.5,29.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_OR2</type>
<position>443,28.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>449.5,28.5</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>413,34</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>412.5,30</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>453,29</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>423,13.5</position>
<gparam>LABEL_TEXT (b) What is the boolean function F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>425.5,-3.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_SMALL_INVERTER</type>
<position>416.5,-2.5</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>406,8.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>406.5,-2.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>406.5,-6.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>402,8.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>400.5,-2.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>401.5,-7</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>453,7</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>445,6.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441,6.5,444,6.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>421.5,7.5,421.5,8.5</points>
<intersection>7.5 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>408,8.5,421.5,8.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>421.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>421.5,7.5,435,7.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>421.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>432,-3.5,432,5.5</points>
<intersection>-3.5 1</intersection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>428.5,-3.5,432,-3.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>432 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>432,5.5,435,5.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>432 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>426.5,31.5,430,31.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>428.5,24.5,430.5,24.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>420,22.5,420,31.5</points>
<intersection>22.5 4</intersection>
<intersection>29.5 2</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>420,31.5,422.5,31.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>420 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>417.5,29.5,420,29.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>420 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>420,22.5,430.5,22.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>420 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>417.5,33.5,430,33.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>417.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>417.5,24.5,417.5,33.5</points>
<intersection>24.5 5</intersection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>417.5,24.5,424.5,24.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>417.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438,29.5,438,32.5</points>
<intersection>29.5 1</intersection>
<intersection>32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>438,29.5,440,29.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>438 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>436,32.5,438,32.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>438 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>438.5,23.5,438.5,27.5</points>
<intersection>23.5 1</intersection>
<intersection>27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>436.5,23.5,438.5,23.5</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>438.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>438.5,27.5,440,27.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>438.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>446,28.5,448.5,28.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<connection>
<GID>52</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>418.5,-2.5,422.5,-2.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>408.5,-2.5,414.5,-2.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>415.5,-6.5,415.5,-4.5</points>
<intersection>-6.5 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>415.5,-4.5,422.5,-4.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>415.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>408.5,-6.5,415.5,-6.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>415.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-37.775,472.076,4.68561,446.463</PageViewport>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>-18,461</position>
<gparam>LABEL_TEXT Design Circuit for F= (A AND (B XOR C)) OR (NOT C)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate></page 6>
<page 7>
<PageViewport>397.9,-83.6854,472.193,-128.501</PageViewport>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>432.5,-103</position>
<gparam>LABEL_TEXT Design Circuit for Truth Table in Ques. - Lecture 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 7>
<page 8>
<PageViewport>878,321.116,1091.21,192.501</PageViewport>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>931.5,303</position>
<gparam>LABEL_TEXT Logic Circuit for overhead light with two switches</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 8>
<page 9>
<PageViewport>997.141,342.896,1916.48,-211.671</PageViewport></page 9></circuit>